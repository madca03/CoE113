`timescale 1ns/1ps
module regfile ( clk, nrst, rd_addrA, rd_addrB, wr_addr, wr_en, wr_data, 
        rd_dataA, rd_dataB );
  input [4:0] rd_addrA;
  input [4:0] rd_addrB;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  output [31:0] rd_dataA;
  output [31:0] rd_dataB;
  input clk, nrst, wr_en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n2000, n2001, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752;
  wire   [31:0] elem01;
  wire   [31:0] elem02;
  wire   [31:0] elem03;
  wire   [31:0] elem04;
  wire   [31:0] elem05;
  wire   [31:0] elem06;
  wire   [31:0] elem07;
  wire   [31:0] elem08;
  wire   [31:0] elem09;
  wire   [31:0] elem10;
  wire   [31:0] elem11;
  wire   [31:0] elem12;
  wire   [31:0] elem13;
  wire   [31:0] elem14;
  wire   [31:0] elem15;
  wire   [31:0] elem16;
  wire   [31:0] elem17;
  wire   [31:0] elem18;
  wire   [31:0] elem19;
  wire   [31:0] elem20;
  wire   [31:0] elem21;
  wire   [31:0] elem22;
  wire   [31:0] elem23;
  wire   [31:0] elem24;
  wire   [31:0] elem25;
  wire   [31:0] elem26;
  wire   [31:0] elem27;
  wire   [31:0] elem28;
  wire   [31:0] elem29;
  wire   [31:0] elem30;
  wire   [31:0] elem31;

  DFFARX1 \elem27_reg[31]  ( .D(n3259), .CLK(clk), .RSTB(n3730), .Q(elem27[31]), .QN(n1) );
  DFFARX1 \elem27_reg[30]  ( .D(n3258), .CLK(clk), .RSTB(n3730), .Q(elem27[30]), .QN(n2) );
  DFFARX1 \elem27_reg[29]  ( .D(n3257), .CLK(clk), .RSTB(n3730), .Q(elem27[29]), .QN(n3) );
  DFFARX1 \elem27_reg[28]  ( .D(n3256), .CLK(clk), .RSTB(n3730), .Q(elem27[28]), .QN(n4) );
  DFFARX1 \elem27_reg[27]  ( .D(n3255), .CLK(clk), .RSTB(n3730), .Q(elem27[27]), .QN(n5) );
  DFFARX1 \elem27_reg[26]  ( .D(n3254), .CLK(clk), .RSTB(n3730), .Q(elem27[26]), .QN(n6) );
  DFFARX1 \elem27_reg[25]  ( .D(n3253), .CLK(clk), .RSTB(n3730), .Q(elem27[25]), .QN(n7) );
  DFFARX1 \elem27_reg[24]  ( .D(n3252), .CLK(clk), .RSTB(n3730), .Q(elem27[24]), .QN(n8) );
  DFFARX1 \elem27_reg[23]  ( .D(n3251), .CLK(clk), .RSTB(n3729), .Q(elem27[23]), .QN(n9) );
  DFFARX1 \elem27_reg[22]  ( .D(n3250), .CLK(clk), .RSTB(n3729), .Q(elem27[22]), .QN(n10) );
  DFFARX1 \elem27_reg[21]  ( .D(n3249), .CLK(clk), .RSTB(n3729), .Q(elem27[21]), .QN(n11) );
  DFFARX1 \elem27_reg[20]  ( .D(n3248), .CLK(clk), .RSTB(n3729), .Q(elem27[20]), .QN(n12) );
  DFFARX1 \elem27_reg[19]  ( .D(n3247), .CLK(clk), .RSTB(n3729), .Q(elem27[19]), .QN(n13) );
  DFFARX1 \elem27_reg[18]  ( .D(n3246), .CLK(clk), .RSTB(n3729), .Q(elem27[18]), .QN(n14) );
  DFFARX1 \elem27_reg[17]  ( .D(n3245), .CLK(clk), .RSTB(n3729), .Q(elem27[17]), .QN(n15) );
  DFFARX1 \elem27_reg[16]  ( .D(n3244), .CLK(clk), .RSTB(n3729), .Q(elem27[16]), .QN(n16) );
  DFFARX1 \elem27_reg[15]  ( .D(n3243), .CLK(clk), .RSTB(n3729), .Q(elem27[15]), .QN(n17) );
  DFFARX1 \elem27_reg[14]  ( .D(n3242), .CLK(clk), .RSTB(n3729), .Q(elem27[14]), .QN(n18) );
  DFFARX1 \elem27_reg[13]  ( .D(n3241), .CLK(clk), .RSTB(n3729), .Q(elem27[13]), .QN(n19) );
  DFFARX1 \elem27_reg[12]  ( .D(n3240), .CLK(clk), .RSTB(n3729), .Q(elem27[12]), .QN(n20) );
  DFFARX1 \elem27_reg[11]  ( .D(n3239), .CLK(clk), .RSTB(n3728), .Q(elem27[11]), .QN(n21) );
  DFFARX1 \elem27_reg[10]  ( .D(n3238), .CLK(clk), .RSTB(n3728), .Q(elem27[10]), .QN(n22) );
  DFFARX1 \elem27_reg[9]  ( .D(n3237), .CLK(clk), .RSTB(n3728), .Q(elem27[9]), 
        .QN(n23) );
  DFFARX1 \elem27_reg[8]  ( .D(n3236), .CLK(clk), .RSTB(n3728), .Q(elem27[8]), 
        .QN(n24) );
  DFFARX1 \elem27_reg[7]  ( .D(n3235), .CLK(clk), .RSTB(n3728), .Q(elem27[7]), 
        .QN(n25) );
  DFFARX1 \elem27_reg[6]  ( .D(n3234), .CLK(clk), .RSTB(n3728), .Q(elem27[6]), 
        .QN(n26) );
  DFFARX1 \elem27_reg[5]  ( .D(n3233), .CLK(clk), .RSTB(n3728), .Q(elem27[5]), 
        .QN(n27) );
  DFFARX1 \elem27_reg[4]  ( .D(n3232), .CLK(clk), .RSTB(n3728), .Q(elem27[4]), 
        .QN(n28) );
  DFFARX1 \elem27_reg[3]  ( .D(n3231), .CLK(clk), .RSTB(n3728), .Q(elem27[3]), 
        .QN(n29) );
  DFFARX1 \elem27_reg[2]  ( .D(n3230), .CLK(clk), .RSTB(n3728), .Q(elem27[2]), 
        .QN(n30) );
  DFFARX1 \elem27_reg[1]  ( .D(n3229), .CLK(clk), .RSTB(n3728), .Q(elem27[1]), 
        .QN(n31) );
  DFFARX1 \elem27_reg[0]  ( .D(n3228), .CLK(clk), .RSTB(n3728), .Q(elem27[0]), 
        .QN(n32) );
  DFFARX1 \elem30_reg[31]  ( .D(n3227), .CLK(clk), .RSTB(n3727), .Q(elem30[31]), .QN(n33) );
  DFFARX1 \elem30_reg[30]  ( .D(n3226), .CLK(clk), .RSTB(n3727), .Q(elem30[30]), .QN(n34) );
  DFFARX1 \elem30_reg[29]  ( .D(n3225), .CLK(clk), .RSTB(n3727), .Q(elem30[29]), .QN(n35) );
  DFFARX1 \elem30_reg[28]  ( .D(n3224), .CLK(clk), .RSTB(n3727), .Q(elem30[28]), .QN(n36) );
  DFFARX1 \elem30_reg[27]  ( .D(n3223), .CLK(clk), .RSTB(n3727), .Q(elem30[27]), .QN(n37) );
  DFFARX1 \elem30_reg[26]  ( .D(n3222), .CLK(clk), .RSTB(n3727), .Q(elem30[26]), .QN(n38) );
  DFFARX1 \elem30_reg[25]  ( .D(n3221), .CLK(clk), .RSTB(n3727), .Q(elem30[25]), .QN(n39) );
  DFFARX1 \elem30_reg[24]  ( .D(n3220), .CLK(clk), .RSTB(n3727), .Q(elem30[24]), .QN(n40) );
  DFFARX1 \elem30_reg[23]  ( .D(n3219), .CLK(clk), .RSTB(n3727), .Q(elem30[23]), .QN(n41) );
  DFFARX1 \elem30_reg[22]  ( .D(n3218), .CLK(clk), .RSTB(n3727), .Q(elem30[22]), .QN(n42) );
  DFFARX1 \elem30_reg[21]  ( .D(n3217), .CLK(clk), .RSTB(n3727), .Q(elem30[21]), .QN(n43) );
  DFFARX1 \elem30_reg[20]  ( .D(n3216), .CLK(clk), .RSTB(n3727), .Q(elem30[20]), .QN(n44) );
  DFFARX1 \elem30_reg[19]  ( .D(n3215), .CLK(clk), .RSTB(n3726), .Q(elem30[19]), .QN(n45) );
  DFFARX1 \elem30_reg[18]  ( .D(n3214), .CLK(clk), .RSTB(n3726), .Q(elem30[18]), .QN(n46) );
  DFFARX1 \elem30_reg[17]  ( .D(n3213), .CLK(clk), .RSTB(n3726), .Q(elem30[17]), .QN(n47) );
  DFFARX1 \elem30_reg[16]  ( .D(n3212), .CLK(clk), .RSTB(n3726), .Q(elem30[16]), .QN(n48) );
  DFFARX1 \elem30_reg[15]  ( .D(n3211), .CLK(clk), .RSTB(n3726), .Q(elem30[15]), .QN(n49) );
  DFFARX1 \elem30_reg[14]  ( .D(n3210), .CLK(clk), .RSTB(n3726), .Q(elem30[14]), .QN(n50) );
  DFFARX1 \elem30_reg[13]  ( .D(n3209), .CLK(clk), .RSTB(n3726), .Q(elem30[13]), .QN(n51) );
  DFFARX1 \elem30_reg[12]  ( .D(n3208), .CLK(clk), .RSTB(n3726), .Q(elem30[12]), .QN(n52) );
  DFFARX1 \elem30_reg[11]  ( .D(n3207), .CLK(clk), .RSTB(n3726), .Q(elem30[11]), .QN(n53) );
  DFFARX1 \elem30_reg[10]  ( .D(n3206), .CLK(clk), .RSTB(n3726), .Q(elem30[10]), .QN(n54) );
  DFFARX1 \elem30_reg[9]  ( .D(n3205), .CLK(clk), .RSTB(n3726), .Q(elem30[9]), 
        .QN(n55) );
  DFFARX1 \elem30_reg[8]  ( .D(n3204), .CLK(clk), .RSTB(n3726), .Q(elem30[8]), 
        .QN(n56) );
  DFFARX1 \elem30_reg[7]  ( .D(n3203), .CLK(clk), .RSTB(n3725), .Q(elem30[7]), 
        .QN(n57) );
  DFFARX1 \elem30_reg[6]  ( .D(n3202), .CLK(clk), .RSTB(n3725), .Q(elem30[6]), 
        .QN(n58) );
  DFFARX1 \elem30_reg[5]  ( .D(n3201), .CLK(clk), .RSTB(n3725), .Q(elem30[5]), 
        .QN(n59) );
  DFFARX1 \elem30_reg[4]  ( .D(n3200), .CLK(clk), .RSTB(n3725), .Q(elem30[4]), 
        .QN(n60) );
  DFFARX1 \elem30_reg[3]  ( .D(n3199), .CLK(clk), .RSTB(n3725), .Q(elem30[3]), 
        .QN(n61) );
  DFFARX1 \elem30_reg[2]  ( .D(n3198), .CLK(clk), .RSTB(n3725), .Q(elem30[2]), 
        .QN(n62) );
  DFFARX1 \elem30_reg[1]  ( .D(n3197), .CLK(clk), .RSTB(n3725), .Q(elem30[1]), 
        .QN(n63) );
  DFFARX1 \elem30_reg[0]  ( .D(n3196), .CLK(clk), .RSTB(n3725), .Q(elem30[0]), 
        .QN(n64) );
  DFFARX1 \elem29_reg[31]  ( .D(n3195), .CLK(clk), .RSTB(n3725), .Q(elem29[31]), .QN(n65) );
  DFFARX1 \elem29_reg[30]  ( .D(n3194), .CLK(clk), .RSTB(n3725), .Q(elem29[30]), .QN(n66) );
  DFFARX1 \elem29_reg[29]  ( .D(n3193), .CLK(clk), .RSTB(n3725), .Q(elem29[29]), .QN(n67) );
  DFFARX1 \elem29_reg[28]  ( .D(n3192), .CLK(clk), .RSTB(n3725), .Q(elem29[28]), .QN(n68) );
  DFFARX1 \elem29_reg[27]  ( .D(n3191), .CLK(clk), .RSTB(n3724), .Q(elem29[27]), .QN(n69) );
  DFFARX1 \elem29_reg[26]  ( .D(n3190), .CLK(clk), .RSTB(n3724), .Q(elem29[26]), .QN(n70) );
  DFFARX1 \elem29_reg[25]  ( .D(n3189), .CLK(clk), .RSTB(n3724), .Q(elem29[25]), .QN(n71) );
  DFFARX1 \elem29_reg[24]  ( .D(n3188), .CLK(clk), .RSTB(n3724), .Q(elem29[24]), .QN(n72) );
  DFFARX1 \elem29_reg[23]  ( .D(n3187), .CLK(clk), .RSTB(n3724), .Q(elem29[23]), .QN(n73) );
  DFFARX1 \elem29_reg[22]  ( .D(n3186), .CLK(clk), .RSTB(n3724), .Q(elem29[22]), .QN(n74) );
  DFFARX1 \elem29_reg[21]  ( .D(n3185), .CLK(clk), .RSTB(n3724), .Q(elem29[21]), .QN(n75) );
  DFFARX1 \elem29_reg[20]  ( .D(n3184), .CLK(clk), .RSTB(n3724), .Q(elem29[20]), .QN(n76) );
  DFFARX1 \elem29_reg[19]  ( .D(n3183), .CLK(clk), .RSTB(n3724), .Q(elem29[19]), .QN(n77) );
  DFFARX1 \elem29_reg[18]  ( .D(n3182), .CLK(clk), .RSTB(n3724), .Q(elem29[18]), .QN(n78) );
  DFFARX1 \elem29_reg[17]  ( .D(n3181), .CLK(clk), .RSTB(n3724), .Q(elem29[17]), .QN(n79) );
  DFFARX1 \elem29_reg[16]  ( .D(n3180), .CLK(clk), .RSTB(n3724), .Q(elem29[16]), .QN(n80) );
  DFFARX1 \elem29_reg[15]  ( .D(n3179), .CLK(clk), .RSTB(n3723), .Q(elem29[15]), .QN(n81) );
  DFFARX1 \elem29_reg[14]  ( .D(n3178), .CLK(clk), .RSTB(n3723), .Q(elem29[14]), .QN(n82) );
  DFFARX1 \elem29_reg[13]  ( .D(n3177), .CLK(clk), .RSTB(n3723), .Q(elem29[13]), .QN(n83) );
  DFFARX1 \elem29_reg[12]  ( .D(n3176), .CLK(clk), .RSTB(n3723), .Q(elem29[12]), .QN(n84) );
  DFFARX1 \elem29_reg[11]  ( .D(n3175), .CLK(clk), .RSTB(n3723), .Q(elem29[11]), .QN(n85) );
  DFFARX1 \elem29_reg[10]  ( .D(n3174), .CLK(clk), .RSTB(n3723), .Q(elem29[10]), .QN(n86) );
  DFFARX1 \elem29_reg[9]  ( .D(n3173), .CLK(clk), .RSTB(n3723), .Q(elem29[9]), 
        .QN(n87) );
  DFFARX1 \elem29_reg[8]  ( .D(n3172), .CLK(clk), .RSTB(n3723), .Q(elem29[8]), 
        .QN(n88) );
  DFFARX1 \elem29_reg[7]  ( .D(n3171), .CLK(clk), .RSTB(n3723), .Q(elem29[7]), 
        .QN(n89) );
  DFFARX1 \elem29_reg[6]  ( .D(n3170), .CLK(clk), .RSTB(n3723), .Q(elem29[6]), 
        .QN(n90) );
  DFFARX1 \elem29_reg[5]  ( .D(n3169), .CLK(clk), .RSTB(n3723), .Q(elem29[5]), 
        .QN(n91) );
  DFFARX1 \elem29_reg[4]  ( .D(n3168), .CLK(clk), .RSTB(n3723), .Q(elem29[4]), 
        .QN(n92) );
  DFFARX1 \elem29_reg[3]  ( .D(n3167), .CLK(clk), .RSTB(n3722), .Q(elem29[3]), 
        .QN(n93) );
  DFFARX1 \elem29_reg[2]  ( .D(n3166), .CLK(clk), .RSTB(n3722), .Q(elem29[2]), 
        .QN(n94) );
  DFFARX1 \elem29_reg[1]  ( .D(n3165), .CLK(clk), .RSTB(n3722), .Q(elem29[1]), 
        .QN(n95) );
  DFFARX1 \elem29_reg[0]  ( .D(n3164), .CLK(clk), .RSTB(n3722), .Q(elem29[0]), 
        .QN(n96) );
  DFFARX1 \elem28_reg[31]  ( .D(n3163), .CLK(clk), .RSTB(n3722), .Q(elem28[31]), .QN(n97) );
  DFFARX1 \elem28_reg[30]  ( .D(n3162), .CLK(clk), .RSTB(n3722), .Q(elem28[30]), .QN(n98) );
  DFFARX1 \elem28_reg[29]  ( .D(n3161), .CLK(clk), .RSTB(n3722), .Q(elem28[29]), .QN(n99) );
  DFFARX1 \elem28_reg[28]  ( .D(n3160), .CLK(clk), .RSTB(n3722), .Q(elem28[28]), .QN(n100) );
  DFFARX1 \elem28_reg[27]  ( .D(n3159), .CLK(clk), .RSTB(n3722), .Q(elem28[27]), .QN(n101) );
  DFFARX1 \elem28_reg[26]  ( .D(n3158), .CLK(clk), .RSTB(n3722), .Q(elem28[26]), .QN(n102) );
  DFFARX1 \elem28_reg[25]  ( .D(n3157), .CLK(clk), .RSTB(n3722), .Q(elem28[25]), .QN(n103) );
  DFFARX1 \elem28_reg[24]  ( .D(n3156), .CLK(clk), .RSTB(n3722), .Q(elem28[24]), .QN(n104) );
  DFFARX1 \elem28_reg[23]  ( .D(n3155), .CLK(clk), .RSTB(n3721), .Q(elem28[23]), .QN(n105) );
  DFFARX1 \elem28_reg[22]  ( .D(n3154), .CLK(clk), .RSTB(n3721), .Q(elem28[22]), .QN(n106) );
  DFFARX1 \elem28_reg[21]  ( .D(n3153), .CLK(clk), .RSTB(n3721), .Q(elem28[21]), .QN(n107) );
  DFFARX1 \elem28_reg[20]  ( .D(n3152), .CLK(clk), .RSTB(n3721), .Q(elem28[20]), .QN(n108) );
  DFFARX1 \elem28_reg[19]  ( .D(n3151), .CLK(clk), .RSTB(n3721), .Q(elem28[19]), .QN(n109) );
  DFFARX1 \elem28_reg[18]  ( .D(n3150), .CLK(clk), .RSTB(n3721), .Q(elem28[18]), .QN(n110) );
  DFFARX1 \elem28_reg[17]  ( .D(n3149), .CLK(clk), .RSTB(n3721), .Q(elem28[17]), .QN(n111) );
  DFFARX1 \elem28_reg[16]  ( .D(n3148), .CLK(clk), .RSTB(n3721), .Q(elem28[16]), .QN(n112) );
  DFFARX1 \elem28_reg[15]  ( .D(n3147), .CLK(clk), .RSTB(n3721), .Q(elem28[15]), .QN(n113) );
  DFFARX1 \elem28_reg[14]  ( .D(n3146), .CLK(clk), .RSTB(n3721), .Q(elem28[14]), .QN(n114) );
  DFFARX1 \elem28_reg[13]  ( .D(n3145), .CLK(clk), .RSTB(n3721), .Q(elem28[13]), .QN(n115) );
  DFFARX1 \elem28_reg[12]  ( .D(n3144), .CLK(clk), .RSTB(n3721), .Q(elem28[12]), .QN(n116) );
  DFFARX1 \elem28_reg[11]  ( .D(n3143), .CLK(clk), .RSTB(n3720), .Q(elem28[11]), .QN(n117) );
  DFFARX1 \elem28_reg[10]  ( .D(n3142), .CLK(clk), .RSTB(n3720), .Q(elem28[10]), .QN(n118) );
  DFFARX1 \elem28_reg[9]  ( .D(n3141), .CLK(clk), .RSTB(n3720), .Q(elem28[9]), 
        .QN(n119) );
  DFFARX1 \elem28_reg[8]  ( .D(n3140), .CLK(clk), .RSTB(n3720), .Q(elem28[8]), 
        .QN(n120) );
  DFFARX1 \elem28_reg[7]  ( .D(n3139), .CLK(clk), .RSTB(n3720), .Q(elem28[7]), 
        .QN(n121) );
  DFFARX1 \elem28_reg[6]  ( .D(n3138), .CLK(clk), .RSTB(n3720), .Q(elem28[6]), 
        .QN(n122) );
  DFFARX1 \elem28_reg[5]  ( .D(n3137), .CLK(clk), .RSTB(n3720), .Q(elem28[5]), 
        .QN(n123) );
  DFFARX1 \elem28_reg[4]  ( .D(n3136), .CLK(clk), .RSTB(n3720), .Q(elem28[4]), 
        .QN(n124) );
  DFFARX1 \elem28_reg[3]  ( .D(n3135), .CLK(clk), .RSTB(n3720), .Q(elem28[3]), 
        .QN(n125) );
  DFFARX1 \elem28_reg[2]  ( .D(n3134), .CLK(clk), .RSTB(n3720), .Q(elem28[2]), 
        .QN(n126) );
  DFFARX1 \elem28_reg[1]  ( .D(n3133), .CLK(clk), .RSTB(n3720), .Q(elem28[1]), 
        .QN(n127) );
  DFFARX1 \elem28_reg[0]  ( .D(n3132), .CLK(clk), .RSTB(n3720), .Q(elem28[0]), 
        .QN(n128) );
  DFFARX1 \elem31_reg[31]  ( .D(n3131), .CLK(clk), .RSTB(n3719), .Q(elem31[31]), .QN(n129) );
  DFFARX1 \elem31_reg[30]  ( .D(n3130), .CLK(clk), .RSTB(n3719), .Q(elem31[30]), .QN(n130) );
  DFFARX1 \elem31_reg[29]  ( .D(n3129), .CLK(clk), .RSTB(n3719), .Q(elem31[29]), .QN(n131) );
  DFFARX1 \elem31_reg[28]  ( .D(n3128), .CLK(clk), .RSTB(n3719), .Q(elem31[28]), .QN(n132) );
  DFFARX1 \elem31_reg[27]  ( .D(n3127), .CLK(clk), .RSTB(n3719), .Q(elem31[27]), .QN(n133) );
  DFFARX1 \elem31_reg[26]  ( .D(n3126), .CLK(clk), .RSTB(n3719), .Q(elem31[26]), .QN(n134) );
  DFFARX1 \elem31_reg[25]  ( .D(n3125), .CLK(clk), .RSTB(n3719), .Q(elem31[25]), .QN(n135) );
  DFFARX1 \elem31_reg[24]  ( .D(n3124), .CLK(clk), .RSTB(n3719), .Q(elem31[24]), .QN(n136) );
  DFFARX1 \elem31_reg[23]  ( .D(n3123), .CLK(clk), .RSTB(n3719), .Q(elem31[23]), .QN(n137) );
  DFFARX1 \elem31_reg[22]  ( .D(n3122), .CLK(clk), .RSTB(n3719), .Q(elem31[22]), .QN(n138) );
  DFFARX1 \elem31_reg[21]  ( .D(n3121), .CLK(clk), .RSTB(n3719), .Q(elem31[21]), .QN(n139) );
  DFFARX1 \elem31_reg[20]  ( .D(n3120), .CLK(clk), .RSTB(n3719), .Q(elem31[20]), .QN(n140) );
  DFFARX1 \elem31_reg[19]  ( .D(n3119), .CLK(clk), .RSTB(n3718), .Q(elem31[19]), .QN(n141) );
  DFFARX1 \elem31_reg[18]  ( .D(n3118), .CLK(clk), .RSTB(n3718), .Q(elem31[18]), .QN(n142) );
  DFFARX1 \elem31_reg[17]  ( .D(n3117), .CLK(clk), .RSTB(n3718), .Q(elem31[17]), .QN(n143) );
  DFFARX1 \elem31_reg[16]  ( .D(n3116), .CLK(clk), .RSTB(n3718), .Q(elem31[16]), .QN(n144) );
  DFFARX1 \elem31_reg[15]  ( .D(n3115), .CLK(clk), .RSTB(n3718), .Q(elem31[15]), .QN(n145) );
  DFFARX1 \elem31_reg[14]  ( .D(n3114), .CLK(clk), .RSTB(n3718), .Q(elem31[14]), .QN(n146) );
  DFFARX1 \elem31_reg[13]  ( .D(n3113), .CLK(clk), .RSTB(n3718), .Q(elem31[13]), .QN(n147) );
  DFFARX1 \elem31_reg[12]  ( .D(n3112), .CLK(clk), .RSTB(n3718), .Q(elem31[12]), .QN(n148) );
  DFFARX1 \elem31_reg[11]  ( .D(n3111), .CLK(clk), .RSTB(n3718), .Q(elem31[11]), .QN(n149) );
  DFFARX1 \elem31_reg[10]  ( .D(n3110), .CLK(clk), .RSTB(n3718), .Q(elem31[10]), .QN(n150) );
  DFFARX1 \elem31_reg[9]  ( .D(n3109), .CLK(clk), .RSTB(n3718), .Q(elem31[9]), 
        .QN(n151) );
  DFFARX1 \elem31_reg[8]  ( .D(n3108), .CLK(clk), .RSTB(n3718), .Q(elem31[8]), 
        .QN(n152) );
  DFFARX1 \elem31_reg[7]  ( .D(n3107), .CLK(clk), .RSTB(n3717), .Q(elem31[7]), 
        .QN(n153) );
  DFFARX1 \elem31_reg[6]  ( .D(n3106), .CLK(clk), .RSTB(n3717), .Q(elem31[6]), 
        .QN(n154) );
  DFFARX1 \elem31_reg[5]  ( .D(n3105), .CLK(clk), .RSTB(n3717), .Q(elem31[5]), 
        .QN(n155) );
  DFFARX1 \elem31_reg[4]  ( .D(n3104), .CLK(clk), .RSTB(n3717), .Q(elem31[4]), 
        .QN(n156) );
  DFFARX1 \elem31_reg[3]  ( .D(n3103), .CLK(clk), .RSTB(n3717), .Q(elem31[3]), 
        .QN(n157) );
  DFFARX1 \elem31_reg[2]  ( .D(n3102), .CLK(clk), .RSTB(n3717), .Q(elem31[2]), 
        .QN(n158) );
  DFFARX1 \elem31_reg[1]  ( .D(n3101), .CLK(clk), .RSTB(n3717), .Q(elem31[1]), 
        .QN(n159) );
  DFFARX1 \elem31_reg[0]  ( .D(n3100), .CLK(clk), .RSTB(n3717), .Q(elem31[0]), 
        .QN(n160) );
  DFFARX1 \elem01_reg[31]  ( .D(n3099), .CLK(clk), .RSTB(n3717), .Q(elem01[31]), .QN(n161) );
  DFFARX1 \elem01_reg[30]  ( .D(n3098), .CLK(clk), .RSTB(n3717), .Q(elem01[30]), .QN(n162) );
  DFFARX1 \elem01_reg[29]  ( .D(n3097), .CLK(clk), .RSTB(n3717), .Q(elem01[29]), .QN(n163) );
  DFFARX1 \elem01_reg[28]  ( .D(n3096), .CLK(clk), .RSTB(n3717), .Q(elem01[28]), .QN(n164) );
  DFFARX1 \elem01_reg[27]  ( .D(n3095), .CLK(clk), .RSTB(n3716), .Q(elem01[27]), .QN(n165) );
  DFFARX1 \elem01_reg[26]  ( .D(n3094), .CLK(clk), .RSTB(n3716), .Q(elem01[26]), .QN(n166) );
  DFFARX1 \elem01_reg[25]  ( .D(n3093), .CLK(clk), .RSTB(n3716), .Q(elem01[25]), .QN(n167) );
  DFFARX1 \elem01_reg[24]  ( .D(n3092), .CLK(clk), .RSTB(n3716), .Q(elem01[24]), .QN(n168) );
  DFFARX1 \elem01_reg[23]  ( .D(n3091), .CLK(clk), .RSTB(n3716), .Q(elem01[23]), .QN(n169) );
  DFFARX1 \elem01_reg[22]  ( .D(n3090), .CLK(clk), .RSTB(n3716), .Q(elem01[22]), .QN(n170) );
  DFFARX1 \elem01_reg[21]  ( .D(n3089), .CLK(clk), .RSTB(n3716), .Q(elem01[21]), .QN(n171) );
  DFFARX1 \elem01_reg[20]  ( .D(n3088), .CLK(clk), .RSTB(n3716), .Q(elem01[20]), .QN(n172) );
  DFFARX1 \elem01_reg[19]  ( .D(n3087), .CLK(clk), .RSTB(n3716), .Q(elem01[19]), .QN(n173) );
  DFFARX1 \elem01_reg[18]  ( .D(n3086), .CLK(clk), .RSTB(n3716), .Q(elem01[18]), .QN(n174) );
  DFFARX1 \elem01_reg[17]  ( .D(n3085), .CLK(clk), .RSTB(n3716), .Q(elem01[17]), .QN(n175) );
  DFFARX1 \elem01_reg[16]  ( .D(n3084), .CLK(clk), .RSTB(n3716), .Q(elem01[16]), .QN(n176) );
  DFFARX1 \elem01_reg[15]  ( .D(n3083), .CLK(clk), .RSTB(n3715), .Q(elem01[15]), .QN(n177) );
  DFFARX1 \elem01_reg[14]  ( .D(n3082), .CLK(clk), .RSTB(n3715), .Q(elem01[14]), .QN(n178) );
  DFFARX1 \elem01_reg[13]  ( .D(n3081), .CLK(clk), .RSTB(n3715), .Q(elem01[13]), .QN(n179) );
  DFFARX1 \elem01_reg[12]  ( .D(n3080), .CLK(clk), .RSTB(n3715), .Q(elem01[12]), .QN(n180) );
  DFFARX1 \elem01_reg[11]  ( .D(n3079), .CLK(clk), .RSTB(n3715), .Q(elem01[11]), .QN(n181) );
  DFFARX1 \elem01_reg[10]  ( .D(n3078), .CLK(clk), .RSTB(n3715), .Q(elem01[10]), .QN(n182) );
  DFFARX1 \elem01_reg[9]  ( .D(n3077), .CLK(clk), .RSTB(n3715), .Q(elem01[9]), 
        .QN(n183) );
  DFFARX1 \elem01_reg[8]  ( .D(n3076), .CLK(clk), .RSTB(n3715), .Q(elem01[8]), 
        .QN(n184) );
  DFFARX1 \elem01_reg[7]  ( .D(n3075), .CLK(clk), .RSTB(n3715), .Q(elem01[7]), 
        .QN(n185) );
  DFFARX1 \elem01_reg[6]  ( .D(n3074), .CLK(clk), .RSTB(n3715), .Q(elem01[6]), 
        .QN(n186) );
  DFFARX1 \elem01_reg[5]  ( .D(n3073), .CLK(clk), .RSTB(n3715), .Q(elem01[5]), 
        .QN(n187) );
  DFFARX1 \elem01_reg[4]  ( .D(n3072), .CLK(clk), .RSTB(n3715), .Q(elem01[4]), 
        .QN(n188) );
  DFFARX1 \elem01_reg[3]  ( .D(n3071), .CLK(clk), .RSTB(n3714), .Q(elem01[3]), 
        .QN(n189) );
  DFFARX1 \elem01_reg[2]  ( .D(n3070), .CLK(clk), .RSTB(n3714), .Q(elem01[2]), 
        .QN(n190) );
  DFFARX1 \elem01_reg[1]  ( .D(n3069), .CLK(clk), .RSTB(n3714), .Q(elem01[1]), 
        .QN(n191) );
  DFFARX1 \elem01_reg[0]  ( .D(n3068), .CLK(clk), .RSTB(n3714), .Q(elem01[0]), 
        .QN(n192) );
  DFFARX1 \elem02_reg[31]  ( .D(n3067), .CLK(clk), .RSTB(n3714), .Q(elem02[31]), .QN(n193) );
  DFFARX1 \elem02_reg[30]  ( .D(n3066), .CLK(clk), .RSTB(n3714), .Q(elem02[30]), .QN(n194) );
  DFFARX1 \elem02_reg[29]  ( .D(n3065), .CLK(clk), .RSTB(n3714), .Q(elem02[29]), .QN(n195) );
  DFFARX1 \elem02_reg[28]  ( .D(n3064), .CLK(clk), .RSTB(n3714), .Q(elem02[28]), .QN(n196) );
  DFFARX1 \elem02_reg[27]  ( .D(n3063), .CLK(clk), .RSTB(n3714), .Q(elem02[27]), .QN(n197) );
  DFFARX1 \elem02_reg[26]  ( .D(n3062), .CLK(clk), .RSTB(n3714), .Q(elem02[26]), .QN(n198) );
  DFFARX1 \elem02_reg[25]  ( .D(n3061), .CLK(clk), .RSTB(n3714), .Q(elem02[25]), .QN(n199) );
  DFFARX1 \elem02_reg[24]  ( .D(n3060), .CLK(clk), .RSTB(n3714), .Q(elem02[24]), .QN(n200) );
  DFFARX1 \elem02_reg[23]  ( .D(n3059), .CLK(clk), .RSTB(n3713), .Q(elem02[23]), .QN(n201) );
  DFFARX1 \elem02_reg[22]  ( .D(n3058), .CLK(clk), .RSTB(n3713), .Q(elem02[22]), .QN(n202) );
  DFFARX1 \elem02_reg[21]  ( .D(n3057), .CLK(clk), .RSTB(n3713), .Q(elem02[21]), .QN(n203) );
  DFFARX1 \elem02_reg[20]  ( .D(n3056), .CLK(clk), .RSTB(n3713), .Q(elem02[20]), .QN(n204) );
  DFFARX1 \elem02_reg[19]  ( .D(n3055), .CLK(clk), .RSTB(n3713), .Q(elem02[19]), .QN(n205) );
  DFFARX1 \elem02_reg[18]  ( .D(n3054), .CLK(clk), .RSTB(n3713), .Q(elem02[18]), .QN(n206) );
  DFFARX1 \elem02_reg[17]  ( .D(n3053), .CLK(clk), .RSTB(n3713), .Q(elem02[17]), .QN(n207) );
  DFFARX1 \elem02_reg[16]  ( .D(n3052), .CLK(clk), .RSTB(n3713), .Q(elem02[16]), .QN(n208) );
  DFFARX1 \elem02_reg[15]  ( .D(n3051), .CLK(clk), .RSTB(n3713), .Q(elem02[15]), .QN(n209) );
  DFFARX1 \elem02_reg[14]  ( .D(n3050), .CLK(clk), .RSTB(n3713), .Q(elem02[14]), .QN(n210) );
  DFFARX1 \elem02_reg[13]  ( .D(n3049), .CLK(clk), .RSTB(n3713), .Q(elem02[13]), .QN(n211) );
  DFFARX1 \elem02_reg[12]  ( .D(n3048), .CLK(clk), .RSTB(n3713), .Q(elem02[12]), .QN(n212) );
  DFFARX1 \elem02_reg[11]  ( .D(n3047), .CLK(clk), .RSTB(n3712), .Q(elem02[11]), .QN(n213) );
  DFFARX1 \elem02_reg[10]  ( .D(n3046), .CLK(clk), .RSTB(n3712), .Q(elem02[10]), .QN(n214) );
  DFFARX1 \elem02_reg[9]  ( .D(n3045), .CLK(clk), .RSTB(n3712), .Q(elem02[9]), 
        .QN(n215) );
  DFFARX1 \elem02_reg[8]  ( .D(n3044), .CLK(clk), .RSTB(n3712), .Q(elem02[8]), 
        .QN(n216) );
  DFFARX1 \elem02_reg[7]  ( .D(n3043), .CLK(clk), .RSTB(n3712), .Q(elem02[7]), 
        .QN(n217) );
  DFFARX1 \elem02_reg[6]  ( .D(n3042), .CLK(clk), .RSTB(n3712), .Q(elem02[6]), 
        .QN(n218) );
  DFFARX1 \elem02_reg[5]  ( .D(n3041), .CLK(clk), .RSTB(n3712), .Q(elem02[5]), 
        .QN(n219) );
  DFFARX1 \elem02_reg[4]  ( .D(n3040), .CLK(clk), .RSTB(n3712), .Q(elem02[4]), 
        .QN(n220) );
  DFFARX1 \elem02_reg[3]  ( .D(n3039), .CLK(clk), .RSTB(n3712), .Q(elem02[3]), 
        .QN(n221) );
  DFFARX1 \elem02_reg[2]  ( .D(n3038), .CLK(clk), .RSTB(n3712), .Q(elem02[2]), 
        .QN(n222) );
  DFFARX1 \elem02_reg[1]  ( .D(n3037), .CLK(clk), .RSTB(n3712), .Q(elem02[1]), 
        .QN(n223) );
  DFFARX1 \elem02_reg[0]  ( .D(n3036), .CLK(clk), .RSTB(n3712), .Q(elem02[0]), 
        .QN(n224) );
  DFFARX1 \elem03_reg[31]  ( .D(n3035), .CLK(clk), .RSTB(n3711), .Q(elem03[31]), .QN(n225) );
  DFFARX1 \elem03_reg[30]  ( .D(n3034), .CLK(clk), .RSTB(n3711), .Q(elem03[30]), .QN(n226) );
  DFFARX1 \elem03_reg[29]  ( .D(n3033), .CLK(clk), .RSTB(n3711), .Q(elem03[29]), .QN(n227) );
  DFFARX1 \elem03_reg[28]  ( .D(n3032), .CLK(clk), .RSTB(n3711), .Q(elem03[28]), .QN(n228) );
  DFFARX1 \elem03_reg[27]  ( .D(n3031), .CLK(clk), .RSTB(n3711), .Q(elem03[27]), .QN(n229) );
  DFFARX1 \elem03_reg[26]  ( .D(n3030), .CLK(clk), .RSTB(n3711), .Q(elem03[26]), .QN(n230) );
  DFFARX1 \elem03_reg[25]  ( .D(n3029), .CLK(clk), .RSTB(n3711), .Q(elem03[25]), .QN(n231) );
  DFFARX1 \elem03_reg[24]  ( .D(n3028), .CLK(clk), .RSTB(n3711), .Q(elem03[24]), .QN(n232) );
  DFFARX1 \elem03_reg[23]  ( .D(n3027), .CLK(clk), .RSTB(n3711), .Q(elem03[23]), .QN(n233) );
  DFFARX1 \elem03_reg[22]  ( .D(n3026), .CLK(clk), .RSTB(n3711), .Q(elem03[22]), .QN(n234) );
  DFFARX1 \elem03_reg[21]  ( .D(n3025), .CLK(clk), .RSTB(n3711), .Q(elem03[21]), .QN(n235) );
  DFFARX1 \elem03_reg[20]  ( .D(n3024), .CLK(clk), .RSTB(n3711), .Q(elem03[20]), .QN(n236) );
  DFFARX1 \elem03_reg[19]  ( .D(n3023), .CLK(clk), .RSTB(n3710), .Q(elem03[19]), .QN(n237) );
  DFFARX1 \elem03_reg[18]  ( .D(n3022), .CLK(clk), .RSTB(n3710), .Q(elem03[18]), .QN(n238) );
  DFFARX1 \elem03_reg[17]  ( .D(n3021), .CLK(clk), .RSTB(n3710), .Q(elem03[17]), .QN(n239) );
  DFFARX1 \elem03_reg[16]  ( .D(n3020), .CLK(clk), .RSTB(n3710), .Q(elem03[16]), .QN(n240) );
  DFFARX1 \elem03_reg[15]  ( .D(n3019), .CLK(clk), .RSTB(n3710), .Q(elem03[15]), .QN(n241) );
  DFFARX1 \elem03_reg[14]  ( .D(n3018), .CLK(clk), .RSTB(n3710), .Q(elem03[14]), .QN(n242) );
  DFFARX1 \elem03_reg[13]  ( .D(n3017), .CLK(clk), .RSTB(n3710), .Q(elem03[13]), .QN(n243) );
  DFFARX1 \elem03_reg[12]  ( .D(n3016), .CLK(clk), .RSTB(n3710), .Q(elem03[12]), .QN(n244) );
  DFFARX1 \elem03_reg[11]  ( .D(n3015), .CLK(clk), .RSTB(n3710), .Q(elem03[11]), .QN(n245) );
  DFFARX1 \elem03_reg[10]  ( .D(n3014), .CLK(clk), .RSTB(n3710), .Q(elem03[10]), .QN(n246) );
  DFFARX1 \elem03_reg[9]  ( .D(n3013), .CLK(clk), .RSTB(n3710), .Q(elem03[9]), 
        .QN(n247) );
  DFFARX1 \elem03_reg[8]  ( .D(n3012), .CLK(clk), .RSTB(n3710), .Q(elem03[8]), 
        .QN(n248) );
  DFFARX1 \elem03_reg[7]  ( .D(n3011), .CLK(clk), .RSTB(n3709), .Q(elem03[7]), 
        .QN(n249) );
  DFFARX1 \elem03_reg[6]  ( .D(n3010), .CLK(clk), .RSTB(n3709), .Q(elem03[6]), 
        .QN(n250) );
  DFFARX1 \elem03_reg[5]  ( .D(n3009), .CLK(clk), .RSTB(n3709), .Q(elem03[5]), 
        .QN(n251) );
  DFFARX1 \elem03_reg[4]  ( .D(n3008), .CLK(clk), .RSTB(n3709), .Q(elem03[4]), 
        .QN(n252) );
  DFFARX1 \elem03_reg[3]  ( .D(n3007), .CLK(clk), .RSTB(n3709), .Q(elem03[3]), 
        .QN(n253) );
  DFFARX1 \elem03_reg[2]  ( .D(n3006), .CLK(clk), .RSTB(n3709), .Q(elem03[2]), 
        .QN(n254) );
  DFFARX1 \elem03_reg[1]  ( .D(n3005), .CLK(clk), .RSTB(n3709), .Q(elem03[1]), 
        .QN(n255) );
  DFFARX1 \elem03_reg[0]  ( .D(n3004), .CLK(clk), .RSTB(n3709), .Q(elem03[0]), 
        .QN(n256) );
  DFFARX1 \elem04_reg[31]  ( .D(n3003), .CLK(clk), .RSTB(n3709), .Q(elem04[31]), .QN(n257) );
  DFFARX1 \elem04_reg[30]  ( .D(n3002), .CLK(clk), .RSTB(n3709), .Q(elem04[30]), .QN(n258) );
  DFFARX1 \elem04_reg[29]  ( .D(n3001), .CLK(clk), .RSTB(n3709), .Q(elem04[29]), .QN(n259) );
  DFFARX1 \elem04_reg[28]  ( .D(n3000), .CLK(clk), .RSTB(n3709), .Q(elem04[28]), .QN(n260) );
  DFFARX1 \elem04_reg[27]  ( .D(n2999), .CLK(clk), .RSTB(n3708), .Q(elem04[27]), .QN(n261) );
  DFFARX1 \elem04_reg[26]  ( .D(n2998), .CLK(clk), .RSTB(n3708), .Q(elem04[26]), .QN(n262) );
  DFFARX1 \elem04_reg[25]  ( .D(n2997), .CLK(clk), .RSTB(n3708), .Q(elem04[25]), .QN(n263) );
  DFFARX1 \elem04_reg[24]  ( .D(n2996), .CLK(clk), .RSTB(n3708), .Q(elem04[24]), .QN(n264) );
  DFFARX1 \elem04_reg[23]  ( .D(n2995), .CLK(clk), .RSTB(n3708), .Q(elem04[23]), .QN(n265) );
  DFFARX1 \elem04_reg[22]  ( .D(n2994), .CLK(clk), .RSTB(n3708), .Q(elem04[22]), .QN(n266) );
  DFFARX1 \elem04_reg[21]  ( .D(n2993), .CLK(clk), .RSTB(n3708), .Q(elem04[21]), .QN(n267) );
  DFFARX1 \elem04_reg[20]  ( .D(n2992), .CLK(clk), .RSTB(n3708), .Q(elem04[20]), .QN(n268) );
  DFFARX1 \elem04_reg[19]  ( .D(n2991), .CLK(clk), .RSTB(n3708), .Q(elem04[19]), .QN(n269) );
  DFFARX1 \elem04_reg[18]  ( .D(n2990), .CLK(clk), .RSTB(n3708), .Q(elem04[18]), .QN(n270) );
  DFFARX1 \elem04_reg[17]  ( .D(n2989), .CLK(clk), .RSTB(n3708), .Q(elem04[17]), .QN(n271) );
  DFFARX1 \elem04_reg[16]  ( .D(n2988), .CLK(clk), .RSTB(n3708), .Q(elem04[16]), .QN(n272) );
  DFFARX1 \elem04_reg[15]  ( .D(n2987), .CLK(clk), .RSTB(n3707), .Q(elem04[15]), .QN(n273) );
  DFFARX1 \elem04_reg[14]  ( .D(n2986), .CLK(clk), .RSTB(n3707), .Q(elem04[14]), .QN(n274) );
  DFFARX1 \elem04_reg[13]  ( .D(n2985), .CLK(clk), .RSTB(n3707), .Q(elem04[13]), .QN(n275) );
  DFFARX1 \elem04_reg[12]  ( .D(n2984), .CLK(clk), .RSTB(n3707), .Q(elem04[12]), .QN(n276) );
  DFFARX1 \elem04_reg[11]  ( .D(n2983), .CLK(clk), .RSTB(n3707), .Q(elem04[11]), .QN(n277) );
  DFFARX1 \elem04_reg[10]  ( .D(n2982), .CLK(clk), .RSTB(n3707), .Q(elem04[10]), .QN(n278) );
  DFFARX1 \elem04_reg[9]  ( .D(n2981), .CLK(clk), .RSTB(n3707), .Q(elem04[9]), 
        .QN(n279) );
  DFFARX1 \elem04_reg[8]  ( .D(n2980), .CLK(clk), .RSTB(n3707), .Q(elem04[8]), 
        .QN(n280) );
  DFFARX1 \elem04_reg[7]  ( .D(n2979), .CLK(clk), .RSTB(n3707), .Q(elem04[7]), 
        .QN(n281) );
  DFFARX1 \elem04_reg[6]  ( .D(n2978), .CLK(clk), .RSTB(n3707), .Q(elem04[6]), 
        .QN(n282) );
  DFFARX1 \elem04_reg[5]  ( .D(n2977), .CLK(clk), .RSTB(n3707), .Q(elem04[5]), 
        .QN(n283) );
  DFFARX1 \elem04_reg[4]  ( .D(n2976), .CLK(clk), .RSTB(n3707), .Q(elem04[4]), 
        .QN(n284) );
  DFFARX1 \elem04_reg[3]  ( .D(n2975), .CLK(clk), .RSTB(n3706), .Q(elem04[3]), 
        .QN(n285) );
  DFFARX1 \elem04_reg[2]  ( .D(n2974), .CLK(clk), .RSTB(n3706), .Q(elem04[2]), 
        .QN(n286) );
  DFFARX1 \elem04_reg[1]  ( .D(n2973), .CLK(clk), .RSTB(n3706), .Q(elem04[1]), 
        .QN(n287) );
  DFFARX1 \elem04_reg[0]  ( .D(n2972), .CLK(clk), .RSTB(n3706), .Q(elem04[0]), 
        .QN(n288) );
  DFFARX1 \elem05_reg[31]  ( .D(n2971), .CLK(clk), .RSTB(n3706), .Q(elem05[31]), .QN(n289) );
  DFFARX1 \elem05_reg[30]  ( .D(n2970), .CLK(clk), .RSTB(n3706), .Q(elem05[30]), .QN(n290) );
  DFFARX1 \elem05_reg[29]  ( .D(n2969), .CLK(clk), .RSTB(n3706), .Q(elem05[29]), .QN(n291) );
  DFFARX1 \elem05_reg[28]  ( .D(n2968), .CLK(clk), .RSTB(n3706), .Q(elem05[28]), .QN(n292) );
  DFFARX1 \elem05_reg[27]  ( .D(n2967), .CLK(clk), .RSTB(n3706), .Q(elem05[27]), .QN(n293) );
  DFFARX1 \elem05_reg[26]  ( .D(n2966), .CLK(clk), .RSTB(n3706), .Q(elem05[26]), .QN(n294) );
  DFFARX1 \elem05_reg[25]  ( .D(n2965), .CLK(clk), .RSTB(n3706), .Q(elem05[25]), .QN(n295) );
  DFFARX1 \elem05_reg[24]  ( .D(n2964), .CLK(clk), .RSTB(n3706), .Q(elem05[24]), .QN(n296) );
  DFFARX1 \elem05_reg[23]  ( .D(n2963), .CLK(clk), .RSTB(n3705), .Q(elem05[23]), .QN(n297) );
  DFFARX1 \elem05_reg[22]  ( .D(n2962), .CLK(clk), .RSTB(n3705), .Q(elem05[22]), .QN(n298) );
  DFFARX1 \elem05_reg[21]  ( .D(n2961), .CLK(clk), .RSTB(n3705), .Q(elem05[21]), .QN(n299) );
  DFFARX1 \elem05_reg[20]  ( .D(n2960), .CLK(clk), .RSTB(n3705), .Q(elem05[20]), .QN(n300) );
  DFFARX1 \elem05_reg[19]  ( .D(n2959), .CLK(clk), .RSTB(n3705), .Q(elem05[19]), .QN(n301) );
  DFFARX1 \elem05_reg[18]  ( .D(n2958), .CLK(clk), .RSTB(n3705), .Q(elem05[18]), .QN(n302) );
  DFFARX1 \elem05_reg[17]  ( .D(n2957), .CLK(clk), .RSTB(n3705), .Q(elem05[17]), .QN(n303) );
  DFFARX1 \elem05_reg[16]  ( .D(n2956), .CLK(clk), .RSTB(n3705), .Q(elem05[16]), .QN(n304) );
  DFFARX1 \elem05_reg[15]  ( .D(n2955), .CLK(clk), .RSTB(n3705), .Q(elem05[15]), .QN(n305) );
  DFFARX1 \elem05_reg[14]  ( .D(n2954), .CLK(clk), .RSTB(n3705), .Q(elem05[14]), .QN(n306) );
  DFFARX1 \elem05_reg[13]  ( .D(n2953), .CLK(clk), .RSTB(n3705), .Q(elem05[13]), .QN(n307) );
  DFFARX1 \elem05_reg[12]  ( .D(n2952), .CLK(clk), .RSTB(n3705), .Q(elem05[12]), .QN(n308) );
  DFFARX1 \elem05_reg[11]  ( .D(n2951), .CLK(clk), .RSTB(n3704), .Q(elem05[11]), .QN(n309) );
  DFFARX1 \elem05_reg[10]  ( .D(n2950), .CLK(clk), .RSTB(n3704), .Q(elem05[10]), .QN(n310) );
  DFFARX1 \elem05_reg[9]  ( .D(n2949), .CLK(clk), .RSTB(n3704), .Q(elem05[9]), 
        .QN(n311) );
  DFFARX1 \elem05_reg[8]  ( .D(n2948), .CLK(clk), .RSTB(n3704), .Q(elem05[8]), 
        .QN(n312) );
  DFFARX1 \elem05_reg[7]  ( .D(n2947), .CLK(clk), .RSTB(n3704), .Q(elem05[7]), 
        .QN(n313) );
  DFFARX1 \elem05_reg[6]  ( .D(n2946), .CLK(clk), .RSTB(n3704), .Q(elem05[6]), 
        .QN(n314) );
  DFFARX1 \elem05_reg[5]  ( .D(n2945), .CLK(clk), .RSTB(n3704), .Q(elem05[5]), 
        .QN(n315) );
  DFFARX1 \elem05_reg[4]  ( .D(n2944), .CLK(clk), .RSTB(n3704), .Q(elem05[4]), 
        .QN(n316) );
  DFFARX1 \elem05_reg[3]  ( .D(n2943), .CLK(clk), .RSTB(n3704), .Q(elem05[3]), 
        .QN(n317) );
  DFFARX1 \elem05_reg[2]  ( .D(n2942), .CLK(clk), .RSTB(n3704), .Q(elem05[2]), 
        .QN(n318) );
  DFFARX1 \elem05_reg[1]  ( .D(n2941), .CLK(clk), .RSTB(n3704), .Q(elem05[1]), 
        .QN(n319) );
  DFFARX1 \elem05_reg[0]  ( .D(n2940), .CLK(clk), .RSTB(n3704), .Q(elem05[0]), 
        .QN(n320) );
  DFFARX1 \elem06_reg[31]  ( .D(n2939), .CLK(clk), .RSTB(n3703), .Q(elem06[31]), .QN(n321) );
  DFFARX1 \elem06_reg[30]  ( .D(n2938), .CLK(clk), .RSTB(n3703), .Q(elem06[30]), .QN(n322) );
  DFFARX1 \elem06_reg[29]  ( .D(n2937), .CLK(clk), .RSTB(n3703), .Q(elem06[29]), .QN(n323) );
  DFFARX1 \elem06_reg[28]  ( .D(n2936), .CLK(clk), .RSTB(n3703), .Q(elem06[28]), .QN(n324) );
  DFFARX1 \elem06_reg[27]  ( .D(n2935), .CLK(clk), .RSTB(n3703), .Q(elem06[27]), .QN(n325) );
  DFFARX1 \elem06_reg[26]  ( .D(n2934), .CLK(clk), .RSTB(n3703), .Q(elem06[26]), .QN(n326) );
  DFFARX1 \elem06_reg[25]  ( .D(n2933), .CLK(clk), .RSTB(n3703), .Q(elem06[25]), .QN(n327) );
  DFFARX1 \elem06_reg[24]  ( .D(n2932), .CLK(clk), .RSTB(n3703), .Q(elem06[24]), .QN(n328) );
  DFFARX1 \elem06_reg[23]  ( .D(n2931), .CLK(clk), .RSTB(n3703), .Q(elem06[23]), .QN(n329) );
  DFFARX1 \elem06_reg[22]  ( .D(n2930), .CLK(clk), .RSTB(n3703), .Q(elem06[22]), .QN(n330) );
  DFFARX1 \elem06_reg[21]  ( .D(n2929), .CLK(clk), .RSTB(n3703), .Q(elem06[21]), .QN(n331) );
  DFFARX1 \elem06_reg[20]  ( .D(n2928), .CLK(clk), .RSTB(n3703), .Q(elem06[20]), .QN(n332) );
  DFFARX1 \elem06_reg[19]  ( .D(n2927), .CLK(clk), .RSTB(n3702), .Q(elem06[19]), .QN(n333) );
  DFFARX1 \elem06_reg[18]  ( .D(n2926), .CLK(clk), .RSTB(n3702), .Q(elem06[18]), .QN(n334) );
  DFFARX1 \elem06_reg[17]  ( .D(n2925), .CLK(clk), .RSTB(n3702), .Q(elem06[17]), .QN(n335) );
  DFFARX1 \elem06_reg[16]  ( .D(n2924), .CLK(clk), .RSTB(n3702), .Q(elem06[16]), .QN(n336) );
  DFFARX1 \elem06_reg[15]  ( .D(n2923), .CLK(clk), .RSTB(n3702), .Q(elem06[15]), .QN(n337) );
  DFFARX1 \elem06_reg[14]  ( .D(n2922), .CLK(clk), .RSTB(n3702), .Q(elem06[14]), .QN(n338) );
  DFFARX1 \elem06_reg[13]  ( .D(n2921), .CLK(clk), .RSTB(n3702), .Q(elem06[13]), .QN(n339) );
  DFFARX1 \elem06_reg[12]  ( .D(n2920), .CLK(clk), .RSTB(n3702), .Q(elem06[12]), .QN(n340) );
  DFFARX1 \elem06_reg[11]  ( .D(n2919), .CLK(clk), .RSTB(n3702), .Q(elem06[11]), .QN(n341) );
  DFFARX1 \elem06_reg[10]  ( .D(n2918), .CLK(clk), .RSTB(n3702), .Q(elem06[10]), .QN(n342) );
  DFFARX1 \elem06_reg[9]  ( .D(n2917), .CLK(clk), .RSTB(n3702), .Q(elem06[9]), 
        .QN(n343) );
  DFFARX1 \elem06_reg[8]  ( .D(n2916), .CLK(clk), .RSTB(n3702), .Q(elem06[8]), 
        .QN(n344) );
  DFFARX1 \elem06_reg[7]  ( .D(n2915), .CLK(clk), .RSTB(n3701), .Q(elem06[7]), 
        .QN(n345) );
  DFFARX1 \elem06_reg[6]  ( .D(n2914), .CLK(clk), .RSTB(n3701), .Q(elem06[6]), 
        .QN(n346) );
  DFFARX1 \elem06_reg[5]  ( .D(n2913), .CLK(clk), .RSTB(n3701), .Q(elem06[5]), 
        .QN(n347) );
  DFFARX1 \elem06_reg[4]  ( .D(n2912), .CLK(clk), .RSTB(n3701), .Q(elem06[4]), 
        .QN(n348) );
  DFFARX1 \elem06_reg[3]  ( .D(n2911), .CLK(clk), .RSTB(n3701), .Q(elem06[3]), 
        .QN(n349) );
  DFFARX1 \elem06_reg[2]  ( .D(n2910), .CLK(clk), .RSTB(n3701), .Q(elem06[2]), 
        .QN(n350) );
  DFFARX1 \elem06_reg[1]  ( .D(n2909), .CLK(clk), .RSTB(n3701), .Q(elem06[1]), 
        .QN(n351) );
  DFFARX1 \elem06_reg[0]  ( .D(n2908), .CLK(clk), .RSTB(n3701), .Q(elem06[0]), 
        .QN(n352) );
  DFFARX1 \elem07_reg[31]  ( .D(n2907), .CLK(clk), .RSTB(n3701), .Q(elem07[31]), .QN(n353) );
  DFFARX1 \elem07_reg[30]  ( .D(n2906), .CLK(clk), .RSTB(n3701), .Q(elem07[30]), .QN(n354) );
  DFFARX1 \elem07_reg[29]  ( .D(n2905), .CLK(clk), .RSTB(n3701), .Q(elem07[29]), .QN(n355) );
  DFFARX1 \elem07_reg[28]  ( .D(n2904), .CLK(clk), .RSTB(n3701), .Q(elem07[28]), .QN(n356) );
  DFFARX1 \elem07_reg[27]  ( .D(n2903), .CLK(clk), .RSTB(n3700), .Q(elem07[27]), .QN(n357) );
  DFFARX1 \elem07_reg[26]  ( .D(n2902), .CLK(clk), .RSTB(n3700), .Q(elem07[26]), .QN(n358) );
  DFFARX1 \elem07_reg[25]  ( .D(n2901), .CLK(clk), .RSTB(n3700), .Q(elem07[25]), .QN(n359) );
  DFFARX1 \elem07_reg[24]  ( .D(n2900), .CLK(clk), .RSTB(n3700), .Q(elem07[24]), .QN(n360) );
  DFFARX1 \elem07_reg[23]  ( .D(n2899), .CLK(clk), .RSTB(n3700), .Q(elem07[23]), .QN(n361) );
  DFFARX1 \elem07_reg[22]  ( .D(n2898), .CLK(clk), .RSTB(n3700), .Q(elem07[22]), .QN(n362) );
  DFFARX1 \elem07_reg[21]  ( .D(n2897), .CLK(clk), .RSTB(n3700), .Q(elem07[21]), .QN(n363) );
  DFFARX1 \elem07_reg[20]  ( .D(n2896), .CLK(clk), .RSTB(n3700), .Q(elem07[20]), .QN(n364) );
  DFFARX1 \elem07_reg[19]  ( .D(n2895), .CLK(clk), .RSTB(n3700), .Q(elem07[19]), .QN(n365) );
  DFFARX1 \elem07_reg[18]  ( .D(n2894), .CLK(clk), .RSTB(n3700), .Q(elem07[18]), .QN(n366) );
  DFFARX1 \elem07_reg[17]  ( .D(n2893), .CLK(clk), .RSTB(n3700), .Q(elem07[17]), .QN(n367) );
  DFFARX1 \elem07_reg[16]  ( .D(n2892), .CLK(clk), .RSTB(n3700), .Q(elem07[16]), .QN(n368) );
  DFFARX1 \elem07_reg[15]  ( .D(n2891), .CLK(clk), .RSTB(n3699), .Q(elem07[15]), .QN(n369) );
  DFFARX1 \elem07_reg[14]  ( .D(n2890), .CLK(clk), .RSTB(n3699), .Q(elem07[14]), .QN(n370) );
  DFFARX1 \elem07_reg[13]  ( .D(n2889), .CLK(clk), .RSTB(n3699), .Q(elem07[13]), .QN(n371) );
  DFFARX1 \elem07_reg[12]  ( .D(n2888), .CLK(clk), .RSTB(n3699), .Q(elem07[12]), .QN(n372) );
  DFFARX1 \elem07_reg[11]  ( .D(n2887), .CLK(clk), .RSTB(n3699), .Q(elem07[11]), .QN(n373) );
  DFFARX1 \elem07_reg[10]  ( .D(n2886), .CLK(clk), .RSTB(n3699), .Q(elem07[10]), .QN(n374) );
  DFFARX1 \elem07_reg[9]  ( .D(n2885), .CLK(clk), .RSTB(n3699), .Q(elem07[9]), 
        .QN(n375) );
  DFFARX1 \elem07_reg[8]  ( .D(n2884), .CLK(clk), .RSTB(n3699), .Q(elem07[8]), 
        .QN(n376) );
  DFFARX1 \elem07_reg[7]  ( .D(n2883), .CLK(clk), .RSTB(n3699), .Q(elem07[7]), 
        .QN(n377) );
  DFFARX1 \elem07_reg[6]  ( .D(n2882), .CLK(clk), .RSTB(n3699), .Q(elem07[6]), 
        .QN(n378) );
  DFFARX1 \elem07_reg[5]  ( .D(n2881), .CLK(clk), .RSTB(n3699), .Q(elem07[5]), 
        .QN(n379) );
  DFFARX1 \elem07_reg[4]  ( .D(n2880), .CLK(clk), .RSTB(n3699), .Q(elem07[4]), 
        .QN(n380) );
  DFFARX1 \elem07_reg[3]  ( .D(n2879), .CLK(clk), .RSTB(n3698), .Q(elem07[3]), 
        .QN(n381) );
  DFFARX1 \elem07_reg[2]  ( .D(n2878), .CLK(clk), .RSTB(n3698), .Q(elem07[2]), 
        .QN(n382) );
  DFFARX1 \elem07_reg[1]  ( .D(n2877), .CLK(clk), .RSTB(n3698), .Q(elem07[1]), 
        .QN(n383) );
  DFFARX1 \elem07_reg[0]  ( .D(n2876), .CLK(clk), .RSTB(n3698), .Q(elem07[0]), 
        .QN(n384) );
  DFFARX1 \elem08_reg[31]  ( .D(n2875), .CLK(clk), .RSTB(n3698), .Q(elem08[31]), .QN(n385) );
  DFFARX1 \elem08_reg[30]  ( .D(n2874), .CLK(clk), .RSTB(n3698), .Q(elem08[30]), .QN(n386) );
  DFFARX1 \elem08_reg[29]  ( .D(n2873), .CLK(clk), .RSTB(n3698), .Q(elem08[29]), .QN(n387) );
  DFFARX1 \elem08_reg[28]  ( .D(n2872), .CLK(clk), .RSTB(n3698), .Q(elem08[28]), .QN(n388) );
  DFFARX1 \elem08_reg[27]  ( .D(n2871), .CLK(clk), .RSTB(n3698), .Q(elem08[27]), .QN(n389) );
  DFFARX1 \elem08_reg[26]  ( .D(n2870), .CLK(clk), .RSTB(n3698), .Q(elem08[26]), .QN(n390) );
  DFFARX1 \elem08_reg[25]  ( .D(n2869), .CLK(clk), .RSTB(n3698), .Q(elem08[25]), .QN(n391) );
  DFFARX1 \elem08_reg[24]  ( .D(n2868), .CLK(clk), .RSTB(n3698), .Q(elem08[24]), .QN(n392) );
  DFFARX1 \elem08_reg[23]  ( .D(n2867), .CLK(clk), .RSTB(n3697), .Q(elem08[23]), .QN(n393) );
  DFFARX1 \elem08_reg[22]  ( .D(n2866), .CLK(clk), .RSTB(n3697), .Q(elem08[22]), .QN(n394) );
  DFFARX1 \elem08_reg[21]  ( .D(n2865), .CLK(clk), .RSTB(n3697), .Q(elem08[21]), .QN(n395) );
  DFFARX1 \elem08_reg[20]  ( .D(n2864), .CLK(clk), .RSTB(n3697), .Q(elem08[20]), .QN(n396) );
  DFFARX1 \elem08_reg[19]  ( .D(n2863), .CLK(clk), .RSTB(n3697), .Q(elem08[19]), .QN(n397) );
  DFFARX1 \elem08_reg[18]  ( .D(n2862), .CLK(clk), .RSTB(n3697), .Q(elem08[18]), .QN(n398) );
  DFFARX1 \elem08_reg[17]  ( .D(n2861), .CLK(clk), .RSTB(n3697), .Q(elem08[17]), .QN(n399) );
  DFFARX1 \elem08_reg[16]  ( .D(n2860), .CLK(clk), .RSTB(n3697), .Q(elem08[16]), .QN(n400) );
  DFFARX1 \elem08_reg[15]  ( .D(n2859), .CLK(clk), .RSTB(n3697), .Q(elem08[15]), .QN(n401) );
  DFFARX1 \elem08_reg[14]  ( .D(n2858), .CLK(clk), .RSTB(n3697), .Q(elem08[14]), .QN(n402) );
  DFFARX1 \elem08_reg[13]  ( .D(n2857), .CLK(clk), .RSTB(n3697), .Q(elem08[13]), .QN(n403) );
  DFFARX1 \elem08_reg[12]  ( .D(n2856), .CLK(clk), .RSTB(n3697), .Q(elem08[12]), .QN(n404) );
  DFFARX1 \elem08_reg[11]  ( .D(n2855), .CLK(clk), .RSTB(n3696), .Q(elem08[11]), .QN(n405) );
  DFFARX1 \elem08_reg[10]  ( .D(n2854), .CLK(clk), .RSTB(n3696), .Q(elem08[10]), .QN(n406) );
  DFFARX1 \elem08_reg[9]  ( .D(n2853), .CLK(clk), .RSTB(n3696), .Q(elem08[9]), 
        .QN(n407) );
  DFFARX1 \elem08_reg[8]  ( .D(n2852), .CLK(clk), .RSTB(n3696), .Q(elem08[8]), 
        .QN(n408) );
  DFFARX1 \elem08_reg[7]  ( .D(n2851), .CLK(clk), .RSTB(n3696), .Q(elem08[7]), 
        .QN(n409) );
  DFFARX1 \elem08_reg[6]  ( .D(n2850), .CLK(clk), .RSTB(n3696), .Q(elem08[6]), 
        .QN(n410) );
  DFFARX1 \elem08_reg[5]  ( .D(n2849), .CLK(clk), .RSTB(n3696), .Q(elem08[5]), 
        .QN(n411) );
  DFFARX1 \elem08_reg[4]  ( .D(n2848), .CLK(clk), .RSTB(n3696), .Q(elem08[4]), 
        .QN(n412) );
  DFFARX1 \elem08_reg[3]  ( .D(n2847), .CLK(clk), .RSTB(n3696), .Q(elem08[3]), 
        .QN(n413) );
  DFFARX1 \elem08_reg[2]  ( .D(n2846), .CLK(clk), .RSTB(n3696), .Q(elem08[2]), 
        .QN(n414) );
  DFFARX1 \elem08_reg[1]  ( .D(n2845), .CLK(clk), .RSTB(n3696), .Q(elem08[1]), 
        .QN(n415) );
  DFFARX1 \elem08_reg[0]  ( .D(n2844), .CLK(clk), .RSTB(n3696), .Q(elem08[0]), 
        .QN(n416) );
  DFFARX1 \elem09_reg[31]  ( .D(n2843), .CLK(clk), .RSTB(n3695), .Q(elem09[31]), .QN(n417) );
  DFFARX1 \elem09_reg[30]  ( .D(n2842), .CLK(clk), .RSTB(n3695), .Q(elem09[30]), .QN(n418) );
  DFFARX1 \elem09_reg[29]  ( .D(n2841), .CLK(clk), .RSTB(n3695), .Q(elem09[29]), .QN(n419) );
  DFFARX1 \elem09_reg[28]  ( .D(n2840), .CLK(clk), .RSTB(n3695), .Q(elem09[28]), .QN(n420) );
  DFFARX1 \elem09_reg[27]  ( .D(n2839), .CLK(clk), .RSTB(n3695), .Q(elem09[27]), .QN(n421) );
  DFFARX1 \elem09_reg[26]  ( .D(n2838), .CLK(clk), .RSTB(n3695), .Q(elem09[26]), .QN(n422) );
  DFFARX1 \elem09_reg[25]  ( .D(n2837), .CLK(clk), .RSTB(n3695), .Q(elem09[25]), .QN(n423) );
  DFFARX1 \elem09_reg[24]  ( .D(n2836), .CLK(clk), .RSTB(n3695), .Q(elem09[24]), .QN(n424) );
  DFFARX1 \elem09_reg[23]  ( .D(n2835), .CLK(clk), .RSTB(n3695), .Q(elem09[23]), .QN(n425) );
  DFFARX1 \elem09_reg[22]  ( .D(n2834), .CLK(clk), .RSTB(n3695), .Q(elem09[22]), .QN(n426) );
  DFFARX1 \elem09_reg[21]  ( .D(n2833), .CLK(clk), .RSTB(n3695), .Q(elem09[21]), .QN(n427) );
  DFFARX1 \elem09_reg[20]  ( .D(n2832), .CLK(clk), .RSTB(n3695), .Q(elem09[20]), .QN(n428) );
  DFFARX1 \elem09_reg[19]  ( .D(n2831), .CLK(clk), .RSTB(n3694), .Q(elem09[19]), .QN(n429) );
  DFFARX1 \elem09_reg[18]  ( .D(n2830), .CLK(clk), .RSTB(n3694), .Q(elem09[18]), .QN(n430) );
  DFFARX1 \elem09_reg[17]  ( .D(n2829), .CLK(clk), .RSTB(n3694), .Q(elem09[17]), .QN(n431) );
  DFFARX1 \elem09_reg[16]  ( .D(n2828), .CLK(clk), .RSTB(n3694), .Q(elem09[16]), .QN(n432) );
  DFFARX1 \elem09_reg[15]  ( .D(n2827), .CLK(clk), .RSTB(n3694), .Q(elem09[15]), .QN(n433) );
  DFFARX1 \elem09_reg[14]  ( .D(n2826), .CLK(clk), .RSTB(n3694), .Q(elem09[14]), .QN(n434) );
  DFFARX1 \elem09_reg[13]  ( .D(n2825), .CLK(clk), .RSTB(n3694), .Q(elem09[13]), .QN(n435) );
  DFFARX1 \elem09_reg[12]  ( .D(n2824), .CLK(clk), .RSTB(n3694), .Q(elem09[12]), .QN(n436) );
  DFFARX1 \elem09_reg[11]  ( .D(n2823), .CLK(clk), .RSTB(n3694), .Q(elem09[11]), .QN(n437) );
  DFFARX1 \elem09_reg[10]  ( .D(n2822), .CLK(clk), .RSTB(n3694), .Q(elem09[10]), .QN(n438) );
  DFFARX1 \elem09_reg[9]  ( .D(n2821), .CLK(clk), .RSTB(n3694), .Q(elem09[9]), 
        .QN(n439) );
  DFFARX1 \elem09_reg[8]  ( .D(n2820), .CLK(clk), .RSTB(n3694), .Q(elem09[8]), 
        .QN(n440) );
  DFFARX1 \elem09_reg[7]  ( .D(n2819), .CLK(clk), .RSTB(n3693), .Q(elem09[7]), 
        .QN(n441) );
  DFFARX1 \elem09_reg[6]  ( .D(n2818), .CLK(clk), .RSTB(n3693), .Q(elem09[6]), 
        .QN(n442) );
  DFFARX1 \elem09_reg[5]  ( .D(n2817), .CLK(clk), .RSTB(n3693), .Q(elem09[5]), 
        .QN(n443) );
  DFFARX1 \elem09_reg[4]  ( .D(n2816), .CLK(clk), .RSTB(n3693), .Q(elem09[4]), 
        .QN(n444) );
  DFFARX1 \elem09_reg[3]  ( .D(n2815), .CLK(clk), .RSTB(n3693), .Q(elem09[3]), 
        .QN(n445) );
  DFFARX1 \elem09_reg[2]  ( .D(n2814), .CLK(clk), .RSTB(n3693), .Q(elem09[2]), 
        .QN(n446) );
  DFFARX1 \elem09_reg[1]  ( .D(n2813), .CLK(clk), .RSTB(n3693), .Q(elem09[1]), 
        .QN(n447) );
  DFFARX1 \elem09_reg[0]  ( .D(n2812), .CLK(clk), .RSTB(n3693), .Q(elem09[0]), 
        .QN(n448) );
  DFFARX1 \elem10_reg[31]  ( .D(n2811), .CLK(clk), .RSTB(n3693), .Q(elem10[31]), .QN(n449) );
  DFFARX1 \elem10_reg[30]  ( .D(n2810), .CLK(clk), .RSTB(n3693), .Q(elem10[30]), .QN(n450) );
  DFFARX1 \elem10_reg[29]  ( .D(n2809), .CLK(clk), .RSTB(n3693), .Q(elem10[29]), .QN(n451) );
  DFFARX1 \elem10_reg[28]  ( .D(n2808), .CLK(clk), .RSTB(n3693), .Q(elem10[28]), .QN(n452) );
  DFFARX1 \elem10_reg[27]  ( .D(n2807), .CLK(clk), .RSTB(n3692), .Q(elem10[27]), .QN(n453) );
  DFFARX1 \elem10_reg[26]  ( .D(n2806), .CLK(clk), .RSTB(n3692), .Q(elem10[26]), .QN(n454) );
  DFFARX1 \elem10_reg[25]  ( .D(n2805), .CLK(clk), .RSTB(n3692), .Q(elem10[25]), .QN(n455) );
  DFFARX1 \elem10_reg[24]  ( .D(n2804), .CLK(clk), .RSTB(n3692), .Q(elem10[24]), .QN(n456) );
  DFFARX1 \elem10_reg[23]  ( .D(n2803), .CLK(clk), .RSTB(n3692), .Q(elem10[23]), .QN(n457) );
  DFFARX1 \elem10_reg[22]  ( .D(n2802), .CLK(clk), .RSTB(n3692), .Q(elem10[22]), .QN(n458) );
  DFFARX1 \elem10_reg[21]  ( .D(n2801), .CLK(clk), .RSTB(n3692), .Q(elem10[21]), .QN(n459) );
  DFFARX1 \elem10_reg[20]  ( .D(n2800), .CLK(clk), .RSTB(n3692), .Q(elem10[20]), .QN(n460) );
  DFFARX1 \elem10_reg[19]  ( .D(n2799), .CLK(clk), .RSTB(n3692), .Q(elem10[19]), .QN(n461) );
  DFFARX1 \elem10_reg[18]  ( .D(n2798), .CLK(clk), .RSTB(n3692), .Q(elem10[18]), .QN(n462) );
  DFFARX1 \elem10_reg[17]  ( .D(n2797), .CLK(clk), .RSTB(n3692), .Q(elem10[17]), .QN(n463) );
  DFFARX1 \elem10_reg[16]  ( .D(n2796), .CLK(clk), .RSTB(n3692), .Q(elem10[16]), .QN(n464) );
  DFFARX1 \elem10_reg[15]  ( .D(n2795), .CLK(clk), .RSTB(n3691), .Q(elem10[15]), .QN(n465) );
  DFFARX1 \elem10_reg[14]  ( .D(n2794), .CLK(clk), .RSTB(n3691), .Q(elem10[14]), .QN(n466) );
  DFFARX1 \elem10_reg[13]  ( .D(n2793), .CLK(clk), .RSTB(n3691), .Q(elem10[13]), .QN(n467) );
  DFFARX1 \elem10_reg[12]  ( .D(n2792), .CLK(clk), .RSTB(n3691), .Q(elem10[12]), .QN(n468) );
  DFFARX1 \elem10_reg[11]  ( .D(n2791), .CLK(clk), .RSTB(n3691), .Q(elem10[11]), .QN(n469) );
  DFFARX1 \elem10_reg[10]  ( .D(n2790), .CLK(clk), .RSTB(n3691), .Q(elem10[10]), .QN(n470) );
  DFFARX1 \elem10_reg[9]  ( .D(n2789), .CLK(clk), .RSTB(n3691), .Q(elem10[9]), 
        .QN(n471) );
  DFFARX1 \elem10_reg[8]  ( .D(n2788), .CLK(clk), .RSTB(n3691), .Q(elem10[8]), 
        .QN(n472) );
  DFFARX1 \elem10_reg[7]  ( .D(n2787), .CLK(clk), .RSTB(n3691), .Q(elem10[7]), 
        .QN(n473) );
  DFFARX1 \elem10_reg[6]  ( .D(n2786), .CLK(clk), .RSTB(n3691), .Q(elem10[6]), 
        .QN(n474) );
  DFFARX1 \elem10_reg[5]  ( .D(n2785), .CLK(clk), .RSTB(n3691), .Q(elem10[5]), 
        .QN(n475) );
  DFFARX1 \elem10_reg[4]  ( .D(n2784), .CLK(clk), .RSTB(n3691), .Q(elem10[4]), 
        .QN(n476) );
  DFFARX1 \elem10_reg[3]  ( .D(n2783), .CLK(clk), .RSTB(n3690), .Q(elem10[3]), 
        .QN(n477) );
  DFFARX1 \elem10_reg[2]  ( .D(n2782), .CLK(clk), .RSTB(n3690), .Q(elem10[2]), 
        .QN(n478) );
  DFFARX1 \elem10_reg[1]  ( .D(n2781), .CLK(clk), .RSTB(n3690), .Q(elem10[1]), 
        .QN(n479) );
  DFFARX1 \elem10_reg[0]  ( .D(n2780), .CLK(clk), .RSTB(n3690), .Q(elem10[0]), 
        .QN(n480) );
  DFFARX1 \elem11_reg[31]  ( .D(n2779), .CLK(clk), .RSTB(n3690), .Q(elem11[31]), .QN(n481) );
  DFFARX1 \elem11_reg[30]  ( .D(n2778), .CLK(clk), .RSTB(n3690), .Q(elem11[30]), .QN(n482) );
  DFFARX1 \elem11_reg[29]  ( .D(n2777), .CLK(clk), .RSTB(n3690), .Q(elem11[29]), .QN(n483) );
  DFFARX1 \elem11_reg[28]  ( .D(n2776), .CLK(clk), .RSTB(n3690), .Q(elem11[28]), .QN(n484) );
  DFFARX1 \elem11_reg[27]  ( .D(n2775), .CLK(clk), .RSTB(n3690), .Q(elem11[27]), .QN(n485) );
  DFFARX1 \elem11_reg[26]  ( .D(n2774), .CLK(clk), .RSTB(n3690), .Q(elem11[26]), .QN(n486) );
  DFFARX1 \elem11_reg[25]  ( .D(n2773), .CLK(clk), .RSTB(n3690), .Q(elem11[25]), .QN(n487) );
  DFFARX1 \elem11_reg[24]  ( .D(n2772), .CLK(clk), .RSTB(n3690), .Q(elem11[24]), .QN(n488) );
  DFFARX1 \elem11_reg[23]  ( .D(n2771), .CLK(clk), .RSTB(n3689), .Q(elem11[23]), .QN(n489) );
  DFFARX1 \elem11_reg[22]  ( .D(n2770), .CLK(clk), .RSTB(n3689), .Q(elem11[22]), .QN(n490) );
  DFFARX1 \elem11_reg[21]  ( .D(n2769), .CLK(clk), .RSTB(n3689), .Q(elem11[21]), .QN(n491) );
  DFFARX1 \elem11_reg[20]  ( .D(n2768), .CLK(clk), .RSTB(n3689), .Q(elem11[20]), .QN(n492) );
  DFFARX1 \elem11_reg[19]  ( .D(n2767), .CLK(clk), .RSTB(n3689), .Q(elem11[19]), .QN(n493) );
  DFFARX1 \elem11_reg[18]  ( .D(n2766), .CLK(clk), .RSTB(n3689), .Q(elem11[18]), .QN(n494) );
  DFFARX1 \elem11_reg[17]  ( .D(n2765), .CLK(clk), .RSTB(n3689), .Q(elem11[17]), .QN(n495) );
  DFFARX1 \elem11_reg[16]  ( .D(n2764), .CLK(clk), .RSTB(n3689), .Q(elem11[16]), .QN(n496) );
  DFFARX1 \elem11_reg[15]  ( .D(n2763), .CLK(clk), .RSTB(n3689), .Q(elem11[15]), .QN(n497) );
  DFFARX1 \elem11_reg[14]  ( .D(n2762), .CLK(clk), .RSTB(n3689), .Q(elem11[14]), .QN(n498) );
  DFFARX1 \elem11_reg[13]  ( .D(n2761), .CLK(clk), .RSTB(n3689), .Q(elem11[13]), .QN(n499) );
  DFFARX1 \elem11_reg[12]  ( .D(n2760), .CLK(clk), .RSTB(n3689), .Q(elem11[12]), .QN(n500) );
  DFFARX1 \elem11_reg[11]  ( .D(n2759), .CLK(clk), .RSTB(n3688), .Q(elem11[11]), .QN(n501) );
  DFFARX1 \elem11_reg[10]  ( .D(n2758), .CLK(clk), .RSTB(n3688), .Q(elem11[10]), .QN(n502) );
  DFFARX1 \elem11_reg[9]  ( .D(n2757), .CLK(clk), .RSTB(n3688), .Q(elem11[9]), 
        .QN(n503) );
  DFFARX1 \elem11_reg[8]  ( .D(n2756), .CLK(clk), .RSTB(n3688), .Q(elem11[8]), 
        .QN(n504) );
  DFFARX1 \elem11_reg[7]  ( .D(n2755), .CLK(clk), .RSTB(n3688), .Q(elem11[7]), 
        .QN(n505) );
  DFFARX1 \elem11_reg[6]  ( .D(n2754), .CLK(clk), .RSTB(n3688), .Q(elem11[6]), 
        .QN(n506) );
  DFFARX1 \elem11_reg[5]  ( .D(n2753), .CLK(clk), .RSTB(n3688), .Q(elem11[5]), 
        .QN(n507) );
  DFFARX1 \elem11_reg[4]  ( .D(n2752), .CLK(clk), .RSTB(n3688), .Q(elem11[4]), 
        .QN(n508) );
  DFFARX1 \elem11_reg[3]  ( .D(n2751), .CLK(clk), .RSTB(n3688), .Q(elem11[3]), 
        .QN(n509) );
  DFFARX1 \elem11_reg[2]  ( .D(n2750), .CLK(clk), .RSTB(n3688), .Q(elem11[2]), 
        .QN(n510) );
  DFFARX1 \elem11_reg[1]  ( .D(n2749), .CLK(clk), .RSTB(n3688), .Q(elem11[1]), 
        .QN(n511) );
  DFFARX1 \elem11_reg[0]  ( .D(n2748), .CLK(clk), .RSTB(n3688), .Q(elem11[0]), 
        .QN(n512) );
  DFFARX1 \elem12_reg[31]  ( .D(n2747), .CLK(clk), .RSTB(n3687), .Q(elem12[31]), .QN(n513) );
  DFFARX1 \elem12_reg[30]  ( .D(n2746), .CLK(clk), .RSTB(n3687), .Q(elem12[30]), .QN(n514) );
  DFFARX1 \elem12_reg[29]  ( .D(n2745), .CLK(clk), .RSTB(n3687), .Q(elem12[29]), .QN(n515) );
  DFFARX1 \elem12_reg[28]  ( .D(n2744), .CLK(clk), .RSTB(n3687), .Q(elem12[28]), .QN(n516) );
  DFFARX1 \elem12_reg[27]  ( .D(n2743), .CLK(clk), .RSTB(n3687), .Q(elem12[27]), .QN(n517) );
  DFFARX1 \elem12_reg[26]  ( .D(n2742), .CLK(clk), .RSTB(n3687), .Q(elem12[26]), .QN(n518) );
  DFFARX1 \elem12_reg[25]  ( .D(n2741), .CLK(clk), .RSTB(n3687), .Q(elem12[25]), .QN(n519) );
  DFFARX1 \elem12_reg[24]  ( .D(n2740), .CLK(clk), .RSTB(n3687), .Q(elem12[24]), .QN(n520) );
  DFFARX1 \elem12_reg[23]  ( .D(n2739), .CLK(clk), .RSTB(n3687), .Q(elem12[23]), .QN(n521) );
  DFFARX1 \elem12_reg[22]  ( .D(n2738), .CLK(clk), .RSTB(n3687), .Q(elem12[22]), .QN(n522) );
  DFFARX1 \elem12_reg[21]  ( .D(n2737), .CLK(clk), .RSTB(n3687), .Q(elem12[21]), .QN(n523) );
  DFFARX1 \elem12_reg[20]  ( .D(n2736), .CLK(clk), .RSTB(n3687), .Q(elem12[20]), .QN(n524) );
  DFFARX1 \elem12_reg[19]  ( .D(n2735), .CLK(clk), .RSTB(n3686), .Q(elem12[19]), .QN(n525) );
  DFFARX1 \elem12_reg[18]  ( .D(n2734), .CLK(clk), .RSTB(n3686), .Q(elem12[18]), .QN(n526) );
  DFFARX1 \elem12_reg[17]  ( .D(n2733), .CLK(clk), .RSTB(n3686), .Q(elem12[17]), .QN(n527) );
  DFFARX1 \elem12_reg[16]  ( .D(n2732), .CLK(clk), .RSTB(n3686), .Q(elem12[16]), .QN(n528) );
  DFFARX1 \elem12_reg[15]  ( .D(n2731), .CLK(clk), .RSTB(n3686), .Q(elem12[15]), .QN(n529) );
  DFFARX1 \elem12_reg[14]  ( .D(n2730), .CLK(clk), .RSTB(n3686), .Q(elem12[14]), .QN(n530) );
  DFFARX1 \elem12_reg[13]  ( .D(n2729), .CLK(clk), .RSTB(n3686), .Q(elem12[13]), .QN(n531) );
  DFFARX1 \elem12_reg[12]  ( .D(n2728), .CLK(clk), .RSTB(n3686), .Q(elem12[12]), .QN(n532) );
  DFFARX1 \elem12_reg[11]  ( .D(n2727), .CLK(clk), .RSTB(n3686), .Q(elem12[11]), .QN(n533) );
  DFFARX1 \elem12_reg[10]  ( .D(n2726), .CLK(clk), .RSTB(n3686), .Q(elem12[10]), .QN(n534) );
  DFFARX1 \elem12_reg[9]  ( .D(n2725), .CLK(clk), .RSTB(n3686), .Q(elem12[9]), 
        .QN(n535) );
  DFFARX1 \elem12_reg[8]  ( .D(n2724), .CLK(clk), .RSTB(n3686), .Q(elem12[8]), 
        .QN(n536) );
  DFFARX1 \elem12_reg[7]  ( .D(n2723), .CLK(clk), .RSTB(n3685), .Q(elem12[7]), 
        .QN(n537) );
  DFFARX1 \elem12_reg[6]  ( .D(n2722), .CLK(clk), .RSTB(n3685), .Q(elem12[6]), 
        .QN(n538) );
  DFFARX1 \elem12_reg[5]  ( .D(n2721), .CLK(clk), .RSTB(n3685), .Q(elem12[5]), 
        .QN(n539) );
  DFFARX1 \elem12_reg[4]  ( .D(n2720), .CLK(clk), .RSTB(n3685), .Q(elem12[4]), 
        .QN(n540) );
  DFFARX1 \elem12_reg[3]  ( .D(n2719), .CLK(clk), .RSTB(n3685), .Q(elem12[3]), 
        .QN(n541) );
  DFFARX1 \elem12_reg[2]  ( .D(n2718), .CLK(clk), .RSTB(n3685), .Q(elem12[2]), 
        .QN(n542) );
  DFFARX1 \elem12_reg[1]  ( .D(n2717), .CLK(clk), .RSTB(n3685), .Q(elem12[1]), 
        .QN(n543) );
  DFFARX1 \elem12_reg[0]  ( .D(n2716), .CLK(clk), .RSTB(n3685), .Q(elem12[0]), 
        .QN(n544) );
  DFFARX1 \elem13_reg[31]  ( .D(n2715), .CLK(clk), .RSTB(n3685), .Q(elem13[31]), .QN(n545) );
  DFFARX1 \elem13_reg[30]  ( .D(n2714), .CLK(clk), .RSTB(n3685), .Q(elem13[30]), .QN(n546) );
  DFFARX1 \elem13_reg[29]  ( .D(n2713), .CLK(clk), .RSTB(n3685), .Q(elem13[29]), .QN(n547) );
  DFFARX1 \elem13_reg[28]  ( .D(n2712), .CLK(clk), .RSTB(n3685), .Q(elem13[28]), .QN(n548) );
  DFFARX1 \elem13_reg[27]  ( .D(n2711), .CLK(clk), .RSTB(n3684), .Q(elem13[27]), .QN(n549) );
  DFFARX1 \elem13_reg[26]  ( .D(n2710), .CLK(clk), .RSTB(n3684), .Q(elem13[26]), .QN(n550) );
  DFFARX1 \elem13_reg[25]  ( .D(n2709), .CLK(clk), .RSTB(n3684), .Q(elem13[25]), .QN(n551) );
  DFFARX1 \elem13_reg[24]  ( .D(n2708), .CLK(clk), .RSTB(n3684), .Q(elem13[24]), .QN(n552) );
  DFFARX1 \elem13_reg[23]  ( .D(n2707), .CLK(clk), .RSTB(n3684), .Q(elem13[23]), .QN(n553) );
  DFFARX1 \elem13_reg[22]  ( .D(n2706), .CLK(clk), .RSTB(n3684), .Q(elem13[22]), .QN(n554) );
  DFFARX1 \elem13_reg[21]  ( .D(n2705), .CLK(clk), .RSTB(n3684), .Q(elem13[21]), .QN(n555) );
  DFFARX1 \elem13_reg[20]  ( .D(n2704), .CLK(clk), .RSTB(n3684), .Q(elem13[20]), .QN(n556) );
  DFFARX1 \elem13_reg[19]  ( .D(n2703), .CLK(clk), .RSTB(n3684), .Q(elem13[19]), .QN(n557) );
  DFFARX1 \elem13_reg[18]  ( .D(n2702), .CLK(clk), .RSTB(n3684), .Q(elem13[18]), .QN(n558) );
  DFFARX1 \elem13_reg[17]  ( .D(n2701), .CLK(clk), .RSTB(n3684), .Q(elem13[17]), .QN(n559) );
  DFFARX1 \elem13_reg[16]  ( .D(n2700), .CLK(clk), .RSTB(n3684), .Q(elem13[16]), .QN(n560) );
  DFFARX1 \elem13_reg[15]  ( .D(n2699), .CLK(clk), .RSTB(n3683), .Q(elem13[15]), .QN(n561) );
  DFFARX1 \elem13_reg[14]  ( .D(n2698), .CLK(clk), .RSTB(n3683), .Q(elem13[14]), .QN(n562) );
  DFFARX1 \elem13_reg[13]  ( .D(n2697), .CLK(clk), .RSTB(n3683), .Q(elem13[13]), .QN(n563) );
  DFFARX1 \elem13_reg[12]  ( .D(n2696), .CLK(clk), .RSTB(n3683), .Q(elem13[12]), .QN(n564) );
  DFFARX1 \elem13_reg[11]  ( .D(n2695), .CLK(clk), .RSTB(n3683), .Q(elem13[11]), .QN(n565) );
  DFFARX1 \elem13_reg[10]  ( .D(n2694), .CLK(clk), .RSTB(n3683), .Q(elem13[10]), .QN(n566) );
  DFFARX1 \elem13_reg[9]  ( .D(n2693), .CLK(clk), .RSTB(n3683), .Q(elem13[9]), 
        .QN(n567) );
  DFFARX1 \elem13_reg[8]  ( .D(n2692), .CLK(clk), .RSTB(n3683), .Q(elem13[8]), 
        .QN(n568) );
  DFFARX1 \elem13_reg[7]  ( .D(n2691), .CLK(clk), .RSTB(n3683), .Q(elem13[7]), 
        .QN(n569) );
  DFFARX1 \elem13_reg[6]  ( .D(n2690), .CLK(clk), .RSTB(n3683), .Q(elem13[6]), 
        .QN(n570) );
  DFFARX1 \elem13_reg[5]  ( .D(n2689), .CLK(clk), .RSTB(n3683), .Q(elem13[5]), 
        .QN(n571) );
  DFFARX1 \elem13_reg[4]  ( .D(n2688), .CLK(clk), .RSTB(n3683), .Q(elem13[4]), 
        .QN(n572) );
  DFFARX1 \elem13_reg[3]  ( .D(n2687), .CLK(clk), .RSTB(n3682), .Q(elem13[3]), 
        .QN(n573) );
  DFFARX1 \elem13_reg[2]  ( .D(n2686), .CLK(clk), .RSTB(n3682), .Q(elem13[2]), 
        .QN(n574) );
  DFFARX1 \elem13_reg[1]  ( .D(n2685), .CLK(clk), .RSTB(n3682), .Q(elem13[1]), 
        .QN(n575) );
  DFFARX1 \elem13_reg[0]  ( .D(n2684), .CLK(clk), .RSTB(n3682), .Q(elem13[0]), 
        .QN(n576) );
  DFFARX1 \elem14_reg[31]  ( .D(n2683), .CLK(clk), .RSTB(n3682), .Q(elem14[31]), .QN(n577) );
  DFFARX1 \elem14_reg[30]  ( .D(n2682), .CLK(clk), .RSTB(n3682), .Q(elem14[30]), .QN(n578) );
  DFFARX1 \elem14_reg[29]  ( .D(n2681), .CLK(clk), .RSTB(n3682), .Q(elem14[29]), .QN(n579) );
  DFFARX1 \elem14_reg[28]  ( .D(n2680), .CLK(clk), .RSTB(n3682), .Q(elem14[28]), .QN(n580) );
  DFFARX1 \elem14_reg[27]  ( .D(n2679), .CLK(clk), .RSTB(n3682), .Q(elem14[27]), .QN(n581) );
  DFFARX1 \elem14_reg[26]  ( .D(n2678), .CLK(clk), .RSTB(n3682), .Q(elem14[26]), .QN(n582) );
  DFFARX1 \elem14_reg[25]  ( .D(n2677), .CLK(clk), .RSTB(n3682), .Q(elem14[25]), .QN(n583) );
  DFFARX1 \elem14_reg[24]  ( .D(n2676), .CLK(clk), .RSTB(n3682), .Q(elem14[24]), .QN(n584) );
  DFFARX1 \elem14_reg[23]  ( .D(n2675), .CLK(clk), .RSTB(n3681), .Q(elem14[23]), .QN(n585) );
  DFFARX1 \elem14_reg[22]  ( .D(n2674), .CLK(clk), .RSTB(n3681), .Q(elem14[22]), .QN(n586) );
  DFFARX1 \elem14_reg[21]  ( .D(n2673), .CLK(clk), .RSTB(n3681), .Q(elem14[21]), .QN(n587) );
  DFFARX1 \elem14_reg[20]  ( .D(n2672), .CLK(clk), .RSTB(n3681), .Q(elem14[20]), .QN(n588) );
  DFFARX1 \elem14_reg[19]  ( .D(n2671), .CLK(clk), .RSTB(n3681), .Q(elem14[19]), .QN(n589) );
  DFFARX1 \elem14_reg[18]  ( .D(n2670), .CLK(clk), .RSTB(n3681), .Q(elem14[18]), .QN(n590) );
  DFFARX1 \elem14_reg[17]  ( .D(n2669), .CLK(clk), .RSTB(n3681), .Q(elem14[17]), .QN(n591) );
  DFFARX1 \elem14_reg[16]  ( .D(n2668), .CLK(clk), .RSTB(n3681), .Q(elem14[16]), .QN(n592) );
  DFFARX1 \elem14_reg[15]  ( .D(n2667), .CLK(clk), .RSTB(n3681), .Q(elem14[15]), .QN(n593) );
  DFFARX1 \elem14_reg[14]  ( .D(n2666), .CLK(clk), .RSTB(n3681), .Q(elem14[14]), .QN(n594) );
  DFFARX1 \elem14_reg[13]  ( .D(n2665), .CLK(clk), .RSTB(n3681), .Q(elem14[13]), .QN(n595) );
  DFFARX1 \elem14_reg[12]  ( .D(n2664), .CLK(clk), .RSTB(n3681), .Q(elem14[12]), .QN(n596) );
  DFFARX1 \elem14_reg[11]  ( .D(n2663), .CLK(clk), .RSTB(n3680), .Q(elem14[11]), .QN(n597) );
  DFFARX1 \elem14_reg[10]  ( .D(n2662), .CLK(clk), .RSTB(n3680), .Q(elem14[10]), .QN(n598) );
  DFFARX1 \elem14_reg[9]  ( .D(n2661), .CLK(clk), .RSTB(n3680), .Q(elem14[9]), 
        .QN(n599) );
  DFFARX1 \elem14_reg[8]  ( .D(n2660), .CLK(clk), .RSTB(n3680), .Q(elem14[8]), 
        .QN(n600) );
  DFFARX1 \elem14_reg[7]  ( .D(n2659), .CLK(clk), .RSTB(n3680), .Q(elem14[7]), 
        .QN(n601) );
  DFFARX1 \elem14_reg[6]  ( .D(n2658), .CLK(clk), .RSTB(n3680), .Q(elem14[6]), 
        .QN(n602) );
  DFFARX1 \elem14_reg[5]  ( .D(n2657), .CLK(clk), .RSTB(n3680), .Q(elem14[5]), 
        .QN(n603) );
  DFFARX1 \elem14_reg[4]  ( .D(n2656), .CLK(clk), .RSTB(n3680), .Q(elem14[4]), 
        .QN(n604) );
  DFFARX1 \elem14_reg[3]  ( .D(n2655), .CLK(clk), .RSTB(n3680), .Q(elem14[3]), 
        .QN(n605) );
  DFFARX1 \elem14_reg[2]  ( .D(n2654), .CLK(clk), .RSTB(n3680), .Q(elem14[2]), 
        .QN(n606) );
  DFFARX1 \elem14_reg[1]  ( .D(n2653), .CLK(clk), .RSTB(n3680), .Q(elem14[1]), 
        .QN(n607) );
  DFFARX1 \elem14_reg[0]  ( .D(n2652), .CLK(clk), .RSTB(n3680), .Q(elem14[0]), 
        .QN(n608) );
  DFFARX1 \elem15_reg[31]  ( .D(n2651), .CLK(clk), .RSTB(n3679), .Q(elem15[31]), .QN(n609) );
  DFFARX1 \elem15_reg[30]  ( .D(n2650), .CLK(clk), .RSTB(n3679), .Q(elem15[30]), .QN(n610) );
  DFFARX1 \elem15_reg[29]  ( .D(n2649), .CLK(clk), .RSTB(n3679), .Q(elem15[29]), .QN(n611) );
  DFFARX1 \elem15_reg[28]  ( .D(n2648), .CLK(clk), .RSTB(n3679), .Q(elem15[28]), .QN(n612) );
  DFFARX1 \elem15_reg[27]  ( .D(n2647), .CLK(clk), .RSTB(n3679), .Q(elem15[27]), .QN(n613) );
  DFFARX1 \elem15_reg[26]  ( .D(n2646), .CLK(clk), .RSTB(n3679), .Q(elem15[26]), .QN(n614) );
  DFFARX1 \elem15_reg[25]  ( .D(n2645), .CLK(clk), .RSTB(n3679), .Q(elem15[25]), .QN(n615) );
  DFFARX1 \elem15_reg[24]  ( .D(n2644), .CLK(clk), .RSTB(n3679), .Q(elem15[24]), .QN(n616) );
  DFFARX1 \elem15_reg[23]  ( .D(n2643), .CLK(clk), .RSTB(n3679), .Q(elem15[23]), .QN(n617) );
  DFFARX1 \elem15_reg[22]  ( .D(n2642), .CLK(clk), .RSTB(n3679), .Q(elem15[22]), .QN(n618) );
  DFFARX1 \elem15_reg[21]  ( .D(n2641), .CLK(clk), .RSTB(n3679), .Q(elem15[21]), .QN(n619) );
  DFFARX1 \elem15_reg[20]  ( .D(n2640), .CLK(clk), .RSTB(n3679), .Q(elem15[20]), .QN(n620) );
  DFFARX1 \elem15_reg[19]  ( .D(n2639), .CLK(clk), .RSTB(n3678), .Q(elem15[19]), .QN(n621) );
  DFFARX1 \elem15_reg[18]  ( .D(n2638), .CLK(clk), .RSTB(n3678), .Q(elem15[18]), .QN(n622) );
  DFFARX1 \elem15_reg[17]  ( .D(n2637), .CLK(clk), .RSTB(n3678), .Q(elem15[17]), .QN(n623) );
  DFFARX1 \elem15_reg[16]  ( .D(n2636), .CLK(clk), .RSTB(n3678), .Q(elem15[16]), .QN(n624) );
  DFFARX1 \elem15_reg[15]  ( .D(n2635), .CLK(clk), .RSTB(n3678), .Q(elem15[15]), .QN(n625) );
  DFFARX1 \elem15_reg[14]  ( .D(n2634), .CLK(clk), .RSTB(n3678), .Q(elem15[14]), .QN(n626) );
  DFFARX1 \elem15_reg[13]  ( .D(n2633), .CLK(clk), .RSTB(n3678), .Q(elem15[13]), .QN(n627) );
  DFFARX1 \elem15_reg[12]  ( .D(n2632), .CLK(clk), .RSTB(n3678), .Q(elem15[12]), .QN(n628) );
  DFFARX1 \elem15_reg[11]  ( .D(n2631), .CLK(clk), .RSTB(n3678), .Q(elem15[11]), .QN(n629) );
  DFFARX1 \elem15_reg[10]  ( .D(n2630), .CLK(clk), .RSTB(n3678), .Q(elem15[10]), .QN(n630) );
  DFFARX1 \elem15_reg[9]  ( .D(n2629), .CLK(clk), .RSTB(n3678), .Q(elem15[9]), 
        .QN(n631) );
  DFFARX1 \elem15_reg[8]  ( .D(n2628), .CLK(clk), .RSTB(n3678), .Q(elem15[8]), 
        .QN(n632) );
  DFFARX1 \elem15_reg[7]  ( .D(n2627), .CLK(clk), .RSTB(n3677), .Q(elem15[7]), 
        .QN(n633) );
  DFFARX1 \elem15_reg[6]  ( .D(n2626), .CLK(clk), .RSTB(n3677), .Q(elem15[6]), 
        .QN(n634) );
  DFFARX1 \elem15_reg[5]  ( .D(n2625), .CLK(clk), .RSTB(n3677), .Q(elem15[5]), 
        .QN(n635) );
  DFFARX1 \elem15_reg[4]  ( .D(n2624), .CLK(clk), .RSTB(n3677), .Q(elem15[4]), 
        .QN(n636) );
  DFFARX1 \elem15_reg[3]  ( .D(n2623), .CLK(clk), .RSTB(n3677), .Q(elem15[3]), 
        .QN(n637) );
  DFFARX1 \elem15_reg[2]  ( .D(n2622), .CLK(clk), .RSTB(n3677), .Q(elem15[2]), 
        .QN(n638) );
  DFFARX1 \elem15_reg[1]  ( .D(n2621), .CLK(clk), .RSTB(n3677), .Q(elem15[1]), 
        .QN(n639) );
  DFFARX1 \elem15_reg[0]  ( .D(n2620), .CLK(clk), .RSTB(n3677), .Q(elem15[0]), 
        .QN(n640) );
  DFFARX1 \elem16_reg[31]  ( .D(n2619), .CLK(clk), .RSTB(n3677), .Q(elem16[31]), .QN(n641) );
  DFFARX1 \elem16_reg[30]  ( .D(n2618), .CLK(clk), .RSTB(n3677), .Q(elem16[30]), .QN(n642) );
  DFFARX1 \elem16_reg[29]  ( .D(n2617), .CLK(clk), .RSTB(n3677), .Q(elem16[29]), .QN(n643) );
  DFFARX1 \elem16_reg[28]  ( .D(n2616), .CLK(clk), .RSTB(n3677), .Q(elem16[28]), .QN(n644) );
  DFFARX1 \elem16_reg[27]  ( .D(n2615), .CLK(clk), .RSTB(n3676), .Q(elem16[27]), .QN(n645) );
  DFFARX1 \elem16_reg[26]  ( .D(n2614), .CLK(clk), .RSTB(n3676), .Q(elem16[26]), .QN(n646) );
  DFFARX1 \elem16_reg[25]  ( .D(n2613), .CLK(clk), .RSTB(n3676), .Q(elem16[25]), .QN(n647) );
  DFFARX1 \elem16_reg[24]  ( .D(n2612), .CLK(clk), .RSTB(n3676), .Q(elem16[24]), .QN(n648) );
  DFFARX1 \elem16_reg[23]  ( .D(n2611), .CLK(clk), .RSTB(n3676), .Q(elem16[23]), .QN(n649) );
  DFFARX1 \elem16_reg[22]  ( .D(n2610), .CLK(clk), .RSTB(n3676), .Q(elem16[22]), .QN(n650) );
  DFFARX1 \elem16_reg[21]  ( .D(n2609), .CLK(clk), .RSTB(n3676), .Q(elem16[21]), .QN(n651) );
  DFFARX1 \elem16_reg[20]  ( .D(n2608), .CLK(clk), .RSTB(n3676), .Q(elem16[20]), .QN(n652) );
  DFFARX1 \elem16_reg[19]  ( .D(n2607), .CLK(clk), .RSTB(n3676), .Q(elem16[19]), .QN(n653) );
  DFFARX1 \elem16_reg[18]  ( .D(n2606), .CLK(clk), .RSTB(n3676), .Q(elem16[18]), .QN(n654) );
  DFFARX1 \elem16_reg[17]  ( .D(n2605), .CLK(clk), .RSTB(n3676), .Q(elem16[17]), .QN(n655) );
  DFFARX1 \elem16_reg[16]  ( .D(n2604), .CLK(clk), .RSTB(n3676), .Q(elem16[16]), .QN(n656) );
  DFFARX1 \elem16_reg[15]  ( .D(n2603), .CLK(clk), .RSTB(n3675), .Q(elem16[15]), .QN(n657) );
  DFFARX1 \elem16_reg[14]  ( .D(n2602), .CLK(clk), .RSTB(n3675), .Q(elem16[14]), .QN(n658) );
  DFFARX1 \elem16_reg[13]  ( .D(n2601), .CLK(clk), .RSTB(n3675), .Q(elem16[13]), .QN(n659) );
  DFFARX1 \elem16_reg[12]  ( .D(n2600), .CLK(clk), .RSTB(n3675), .Q(elem16[12]), .QN(n660) );
  DFFARX1 \elem16_reg[11]  ( .D(n2599), .CLK(clk), .RSTB(n3675), .Q(elem16[11]), .QN(n661) );
  DFFARX1 \elem16_reg[10]  ( .D(n2598), .CLK(clk), .RSTB(n3675), .Q(elem16[10]), .QN(n662) );
  DFFARX1 \elem16_reg[9]  ( .D(n2597), .CLK(clk), .RSTB(n3675), .Q(elem16[9]), 
        .QN(n663) );
  DFFARX1 \elem16_reg[8]  ( .D(n2596), .CLK(clk), .RSTB(n3675), .Q(elem16[8]), 
        .QN(n664) );
  DFFARX1 \elem16_reg[7]  ( .D(n2595), .CLK(clk), .RSTB(n3675), .Q(elem16[7]), 
        .QN(n665) );
  DFFARX1 \elem16_reg[6]  ( .D(n2594), .CLK(clk), .RSTB(n3675), .Q(elem16[6]), 
        .QN(n666) );
  DFFARX1 \elem16_reg[5]  ( .D(n2593), .CLK(clk), .RSTB(n3675), .Q(elem16[5]), 
        .QN(n667) );
  DFFARX1 \elem16_reg[4]  ( .D(n2592), .CLK(clk), .RSTB(n3675), .Q(elem16[4]), 
        .QN(n668) );
  DFFARX1 \elem16_reg[3]  ( .D(n2591), .CLK(clk), .RSTB(n3674), .Q(elem16[3]), 
        .QN(n669) );
  DFFARX1 \elem16_reg[2]  ( .D(n2590), .CLK(clk), .RSTB(n3674), .Q(elem16[2]), 
        .QN(n670) );
  DFFARX1 \elem16_reg[1]  ( .D(n2589), .CLK(clk), .RSTB(n3674), .Q(elem16[1]), 
        .QN(n671) );
  DFFARX1 \elem16_reg[0]  ( .D(n2588), .CLK(clk), .RSTB(n3674), .Q(elem16[0]), 
        .QN(n672) );
  DFFARX1 \elem17_reg[31]  ( .D(n2587), .CLK(clk), .RSTB(n3674), .Q(elem17[31]), .QN(n673) );
  DFFARX1 \elem17_reg[30]  ( .D(n2586), .CLK(clk), .RSTB(n3674), .Q(elem17[30]), .QN(n674) );
  DFFARX1 \elem17_reg[29]  ( .D(n2585), .CLK(clk), .RSTB(n3674), .Q(elem17[29]), .QN(n675) );
  DFFARX1 \elem17_reg[28]  ( .D(n2584), .CLK(clk), .RSTB(n3674), .Q(elem17[28]), .QN(n676) );
  DFFARX1 \elem17_reg[27]  ( .D(n2583), .CLK(clk), .RSTB(n3674), .Q(elem17[27]), .QN(n677) );
  DFFARX1 \elem17_reg[26]  ( .D(n2582), .CLK(clk), .RSTB(n3674), .Q(elem17[26]), .QN(n678) );
  DFFARX1 \elem17_reg[25]  ( .D(n2581), .CLK(clk), .RSTB(n3674), .Q(elem17[25]), .QN(n679) );
  DFFARX1 \elem17_reg[24]  ( .D(n2580), .CLK(clk), .RSTB(n3674), .Q(elem17[24]), .QN(n680) );
  DFFARX1 \elem17_reg[23]  ( .D(n2579), .CLK(clk), .RSTB(n3673), .Q(elem17[23]), .QN(n681) );
  DFFARX1 \elem17_reg[22]  ( .D(n2578), .CLK(clk), .RSTB(n3673), .Q(elem17[22]), .QN(n682) );
  DFFARX1 \elem17_reg[21]  ( .D(n2577), .CLK(clk), .RSTB(n3673), .Q(elem17[21]), .QN(n683) );
  DFFARX1 \elem17_reg[20]  ( .D(n2576), .CLK(clk), .RSTB(n3673), .Q(elem17[20]), .QN(n684) );
  DFFARX1 \elem17_reg[19]  ( .D(n2575), .CLK(clk), .RSTB(n3673), .Q(elem17[19]), .QN(n685) );
  DFFARX1 \elem17_reg[18]  ( .D(n2574), .CLK(clk), .RSTB(n3673), .Q(elem17[18]), .QN(n686) );
  DFFARX1 \elem17_reg[17]  ( .D(n2573), .CLK(clk), .RSTB(n3673), .Q(elem17[17]), .QN(n687) );
  DFFARX1 \elem17_reg[16]  ( .D(n2572), .CLK(clk), .RSTB(n3673), .Q(elem17[16]), .QN(n688) );
  DFFARX1 \elem17_reg[15]  ( .D(n2571), .CLK(clk), .RSTB(n3673), .Q(elem17[15]), .QN(n689) );
  DFFARX1 \elem17_reg[14]  ( .D(n2570), .CLK(clk), .RSTB(n3673), .Q(elem17[14]), .QN(n690) );
  DFFARX1 \elem17_reg[13]  ( .D(n2569), .CLK(clk), .RSTB(n3673), .Q(elem17[13]), .QN(n691) );
  DFFARX1 \elem17_reg[12]  ( .D(n2568), .CLK(clk), .RSTB(n3673), .Q(elem17[12]), .QN(n692) );
  DFFARX1 \elem17_reg[11]  ( .D(n2567), .CLK(clk), .RSTB(n3672), .Q(elem17[11]), .QN(n693) );
  DFFARX1 \elem17_reg[10]  ( .D(n2566), .CLK(clk), .RSTB(n3672), .Q(elem17[10]), .QN(n694) );
  DFFARX1 \elem17_reg[9]  ( .D(n2565), .CLK(clk), .RSTB(n3672), .Q(elem17[9]), 
        .QN(n695) );
  DFFARX1 \elem17_reg[8]  ( .D(n2564), .CLK(clk), .RSTB(n3672), .Q(elem17[8]), 
        .QN(n696) );
  DFFARX1 \elem17_reg[7]  ( .D(n2563), .CLK(clk), .RSTB(n3672), .Q(elem17[7]), 
        .QN(n697) );
  DFFARX1 \elem17_reg[6]  ( .D(n2562), .CLK(clk), .RSTB(n3672), .Q(elem17[6]), 
        .QN(n698) );
  DFFARX1 \elem17_reg[5]  ( .D(n2561), .CLK(clk), .RSTB(n3672), .Q(elem17[5]), 
        .QN(n699) );
  DFFARX1 \elem17_reg[4]  ( .D(n2560), .CLK(clk), .RSTB(n3672), .Q(elem17[4]), 
        .QN(n700) );
  DFFARX1 \elem17_reg[3]  ( .D(n2559), .CLK(clk), .RSTB(n3672), .Q(elem17[3]), 
        .QN(n701) );
  DFFARX1 \elem17_reg[2]  ( .D(n2558), .CLK(clk), .RSTB(n3672), .Q(elem17[2]), 
        .QN(n702) );
  DFFARX1 \elem17_reg[1]  ( .D(n2557), .CLK(clk), .RSTB(n3672), .Q(elem17[1]), 
        .QN(n703) );
  DFFARX1 \elem17_reg[0]  ( .D(n2556), .CLK(clk), .RSTB(n3672), .Q(elem17[0]), 
        .QN(n704) );
  DFFARX1 \elem18_reg[31]  ( .D(n2555), .CLK(clk), .RSTB(n3671), .Q(elem18[31]), .QN(n705) );
  DFFARX1 \elem18_reg[30]  ( .D(n2554), .CLK(clk), .RSTB(n3671), .Q(elem18[30]), .QN(n706) );
  DFFARX1 \elem18_reg[29]  ( .D(n2553), .CLK(clk), .RSTB(n3671), .Q(elem18[29]), .QN(n707) );
  DFFARX1 \elem18_reg[28]  ( .D(n2552), .CLK(clk), .RSTB(n3671), .Q(elem18[28]), .QN(n708) );
  DFFARX1 \elem18_reg[27]  ( .D(n2551), .CLK(clk), .RSTB(n3671), .Q(elem18[27]), .QN(n709) );
  DFFARX1 \elem18_reg[26]  ( .D(n2550), .CLK(clk), .RSTB(n3671), .Q(elem18[26]), .QN(n710) );
  DFFARX1 \elem18_reg[25]  ( .D(n2549), .CLK(clk), .RSTB(n3671), .Q(elem18[25]), .QN(n711) );
  DFFARX1 \elem18_reg[24]  ( .D(n2548), .CLK(clk), .RSTB(n3671), .Q(elem18[24]), .QN(n712) );
  DFFARX1 \elem18_reg[23]  ( .D(n2547), .CLK(clk), .RSTB(n3671), .Q(elem18[23]), .QN(n713) );
  DFFARX1 \elem18_reg[22]  ( .D(n2546), .CLK(clk), .RSTB(n3671), .Q(elem18[22]), .QN(n714) );
  DFFARX1 \elem18_reg[21]  ( .D(n2545), .CLK(clk), .RSTB(n3671), .Q(elem18[21]), .QN(n715) );
  DFFARX1 \elem18_reg[20]  ( .D(n2544), .CLK(clk), .RSTB(n3671), .Q(elem18[20]), .QN(n716) );
  DFFARX1 \elem18_reg[19]  ( .D(n2543), .CLK(clk), .RSTB(n3670), .Q(elem18[19]), .QN(n717) );
  DFFARX1 \elem18_reg[18]  ( .D(n2542), .CLK(clk), .RSTB(n3670), .Q(elem18[18]), .QN(n718) );
  DFFARX1 \elem18_reg[17]  ( .D(n2541), .CLK(clk), .RSTB(n3670), .Q(elem18[17]), .QN(n719) );
  DFFARX1 \elem18_reg[16]  ( .D(n2540), .CLK(clk), .RSTB(n3670), .Q(elem18[16]), .QN(n720) );
  DFFARX1 \elem18_reg[15]  ( .D(n2539), .CLK(clk), .RSTB(n3670), .Q(elem18[15]), .QN(n721) );
  DFFARX1 \elem18_reg[14]  ( .D(n2538), .CLK(clk), .RSTB(n3670), .Q(elem18[14]), .QN(n722) );
  DFFARX1 \elem18_reg[13]  ( .D(n2537), .CLK(clk), .RSTB(n3670), .Q(elem18[13]), .QN(n723) );
  DFFARX1 \elem18_reg[12]  ( .D(n2536), .CLK(clk), .RSTB(n3670), .Q(elem18[12]), .QN(n724) );
  DFFARX1 \elem18_reg[11]  ( .D(n2535), .CLK(clk), .RSTB(n3670), .Q(elem18[11]), .QN(n725) );
  DFFARX1 \elem18_reg[10]  ( .D(n2534), .CLK(clk), .RSTB(n3670), .Q(elem18[10]), .QN(n726) );
  DFFARX1 \elem18_reg[9]  ( .D(n2533), .CLK(clk), .RSTB(n3670), .Q(elem18[9]), 
        .QN(n727) );
  DFFARX1 \elem18_reg[8]  ( .D(n2532), .CLK(clk), .RSTB(n3670), .Q(elem18[8]), 
        .QN(n728) );
  DFFARX1 \elem18_reg[7]  ( .D(n2531), .CLK(clk), .RSTB(n3669), .Q(elem18[7]), 
        .QN(n729) );
  DFFARX1 \elem18_reg[6]  ( .D(n2530), .CLK(clk), .RSTB(n3669), .Q(elem18[6]), 
        .QN(n730) );
  DFFARX1 \elem18_reg[5]  ( .D(n2529), .CLK(clk), .RSTB(n3669), .Q(elem18[5]), 
        .QN(n731) );
  DFFARX1 \elem18_reg[4]  ( .D(n2528), .CLK(clk), .RSTB(n3669), .Q(elem18[4]), 
        .QN(n732) );
  DFFARX1 \elem18_reg[3]  ( .D(n2527), .CLK(clk), .RSTB(n3669), .Q(elem18[3]), 
        .QN(n733) );
  DFFARX1 \elem18_reg[2]  ( .D(n2526), .CLK(clk), .RSTB(n3669), .Q(elem18[2]), 
        .QN(n734) );
  DFFARX1 \elem18_reg[1]  ( .D(n2525), .CLK(clk), .RSTB(n3669), .Q(elem18[1]), 
        .QN(n735) );
  DFFARX1 \elem18_reg[0]  ( .D(n2524), .CLK(clk), .RSTB(n3669), .Q(elem18[0]), 
        .QN(n736) );
  DFFARX1 \elem19_reg[31]  ( .D(n2523), .CLK(clk), .RSTB(n3669), .Q(elem19[31]), .QN(n737) );
  DFFARX1 \elem19_reg[30]  ( .D(n2522), .CLK(clk), .RSTB(n3669), .Q(elem19[30]), .QN(n738) );
  DFFARX1 \elem19_reg[29]  ( .D(n2521), .CLK(clk), .RSTB(n3669), .Q(elem19[29]), .QN(n739) );
  DFFARX1 \elem19_reg[28]  ( .D(n2520), .CLK(clk), .RSTB(n3669), .Q(elem19[28]), .QN(n740) );
  DFFARX1 \elem19_reg[27]  ( .D(n2519), .CLK(clk), .RSTB(n3668), .Q(elem19[27]), .QN(n741) );
  DFFARX1 \elem19_reg[26]  ( .D(n2518), .CLK(clk), .RSTB(n3668), .Q(elem19[26]), .QN(n742) );
  DFFARX1 \elem19_reg[25]  ( .D(n2517), .CLK(clk), .RSTB(n3668), .Q(elem19[25]), .QN(n743) );
  DFFARX1 \elem19_reg[24]  ( .D(n2516), .CLK(clk), .RSTB(n3668), .Q(elem19[24]), .QN(n744) );
  DFFARX1 \elem19_reg[23]  ( .D(n2515), .CLK(clk), .RSTB(n3668), .Q(elem19[23]), .QN(n745) );
  DFFARX1 \elem19_reg[22]  ( .D(n2514), .CLK(clk), .RSTB(n3668), .Q(elem19[22]), .QN(n746) );
  DFFARX1 \elem19_reg[21]  ( .D(n2513), .CLK(clk), .RSTB(n3668), .Q(elem19[21]), .QN(n747) );
  DFFARX1 \elem19_reg[20]  ( .D(n2512), .CLK(clk), .RSTB(n3668), .Q(elem19[20]), .QN(n748) );
  DFFARX1 \elem19_reg[19]  ( .D(n2511), .CLK(clk), .RSTB(n3668), .Q(elem19[19]), .QN(n749) );
  DFFARX1 \elem19_reg[18]  ( .D(n2510), .CLK(clk), .RSTB(n3668), .Q(elem19[18]), .QN(n750) );
  DFFARX1 \elem19_reg[17]  ( .D(n2509), .CLK(clk), .RSTB(n3668), .Q(elem19[17]), .QN(n751) );
  DFFARX1 \elem19_reg[16]  ( .D(n2508), .CLK(clk), .RSTB(n3668), .Q(elem19[16]), .QN(n752) );
  DFFARX1 \elem19_reg[15]  ( .D(n2507), .CLK(clk), .RSTB(n3667), .Q(elem19[15]), .QN(n753) );
  DFFARX1 \elem19_reg[14]  ( .D(n2506), .CLK(clk), .RSTB(n3667), .Q(elem19[14]), .QN(n754) );
  DFFARX1 \elem19_reg[13]  ( .D(n2505), .CLK(clk), .RSTB(n3667), .Q(elem19[13]), .QN(n755) );
  DFFARX1 \elem19_reg[12]  ( .D(n2504), .CLK(clk), .RSTB(n3667), .Q(elem19[12]), .QN(n756) );
  DFFARX1 \elem19_reg[11]  ( .D(n2503), .CLK(clk), .RSTB(n3667), .Q(elem19[11]), .QN(n757) );
  DFFARX1 \elem19_reg[10]  ( .D(n2502), .CLK(clk), .RSTB(n3667), .Q(elem19[10]), .QN(n758) );
  DFFARX1 \elem19_reg[9]  ( .D(n2501), .CLK(clk), .RSTB(n3667), .Q(elem19[9]), 
        .QN(n759) );
  DFFARX1 \elem19_reg[8]  ( .D(n2500), .CLK(clk), .RSTB(n3667), .Q(elem19[8]), 
        .QN(n760) );
  DFFARX1 \elem19_reg[7]  ( .D(n2499), .CLK(clk), .RSTB(n3667), .Q(elem19[7]), 
        .QN(n761) );
  DFFARX1 \elem19_reg[6]  ( .D(n2498), .CLK(clk), .RSTB(n3667), .Q(elem19[6]), 
        .QN(n762) );
  DFFARX1 \elem19_reg[5]  ( .D(n2497), .CLK(clk), .RSTB(n3667), .Q(elem19[5]), 
        .QN(n763) );
  DFFARX1 \elem19_reg[4]  ( .D(n2496), .CLK(clk), .RSTB(n3667), .Q(elem19[4]), 
        .QN(n764) );
  DFFARX1 \elem19_reg[3]  ( .D(n2495), .CLK(clk), .RSTB(n3666), .Q(elem19[3]), 
        .QN(n765) );
  DFFARX1 \elem19_reg[2]  ( .D(n2494), .CLK(clk), .RSTB(n3666), .Q(elem19[2]), 
        .QN(n766) );
  DFFARX1 \elem19_reg[1]  ( .D(n2493), .CLK(clk), .RSTB(n3666), .Q(elem19[1]), 
        .QN(n767) );
  DFFARX1 \elem19_reg[0]  ( .D(n2492), .CLK(clk), .RSTB(n3666), .Q(elem19[0]), 
        .QN(n768) );
  DFFARX1 \elem20_reg[31]  ( .D(n2491), .CLK(clk), .RSTB(n3666), .Q(elem20[31]), .QN(n769) );
  DFFARX1 \elem20_reg[30]  ( .D(n2490), .CLK(clk), .RSTB(n3666), .Q(elem20[30]), .QN(n770) );
  DFFARX1 \elem20_reg[29]  ( .D(n2489), .CLK(clk), .RSTB(n3666), .Q(elem20[29]), .QN(n771) );
  DFFARX1 \elem20_reg[28]  ( .D(n2488), .CLK(clk), .RSTB(n3666), .Q(elem20[28]), .QN(n772) );
  DFFARX1 \elem20_reg[27]  ( .D(n2487), .CLK(clk), .RSTB(n3666), .Q(elem20[27]), .QN(n773) );
  DFFARX1 \elem20_reg[26]  ( .D(n2486), .CLK(clk), .RSTB(n3666), .Q(elem20[26]), .QN(n774) );
  DFFARX1 \elem20_reg[25]  ( .D(n2485), .CLK(clk), .RSTB(n3666), .Q(elem20[25]), .QN(n775) );
  DFFARX1 \elem20_reg[24]  ( .D(n2484), .CLK(clk), .RSTB(n3666), .Q(elem20[24]), .QN(n776) );
  DFFARX1 \elem20_reg[23]  ( .D(n2483), .CLK(clk), .RSTB(n3665), .Q(elem20[23]), .QN(n777) );
  DFFARX1 \elem20_reg[22]  ( .D(n2482), .CLK(clk), .RSTB(n3665), .Q(elem20[22]), .QN(n778) );
  DFFARX1 \elem20_reg[21]  ( .D(n2481), .CLK(clk), .RSTB(n3665), .Q(elem20[21]), .QN(n779) );
  DFFARX1 \elem20_reg[20]  ( .D(n2480), .CLK(clk), .RSTB(n3665), .Q(elem20[20]), .QN(n780) );
  DFFARX1 \elem20_reg[19]  ( .D(n2479), .CLK(clk), .RSTB(n3665), .Q(elem20[19]), .QN(n781) );
  DFFARX1 \elem20_reg[18]  ( .D(n2478), .CLK(clk), .RSTB(n3665), .Q(elem20[18]), .QN(n782) );
  DFFARX1 \elem20_reg[17]  ( .D(n2477), .CLK(clk), .RSTB(n3665), .Q(elem20[17]), .QN(n783) );
  DFFARX1 \elem20_reg[16]  ( .D(n2476), .CLK(clk), .RSTB(n3665), .Q(elem20[16]), .QN(n784) );
  DFFARX1 \elem20_reg[15]  ( .D(n2475), .CLK(clk), .RSTB(n3665), .Q(elem20[15]), .QN(n785) );
  DFFARX1 \elem20_reg[14]  ( .D(n2474), .CLK(clk), .RSTB(n3665), .Q(elem20[14]), .QN(n786) );
  DFFARX1 \elem20_reg[13]  ( .D(n2473), .CLK(clk), .RSTB(n3665), .Q(elem20[13]), .QN(n787) );
  DFFARX1 \elem20_reg[12]  ( .D(n2472), .CLK(clk), .RSTB(n3665), .Q(elem20[12]), .QN(n788) );
  DFFARX1 \elem20_reg[11]  ( .D(n2471), .CLK(clk), .RSTB(n3664), .Q(elem20[11]), .QN(n789) );
  DFFARX1 \elem20_reg[10]  ( .D(n2470), .CLK(clk), .RSTB(n3664), .Q(elem20[10]), .QN(n790) );
  DFFARX1 \elem20_reg[9]  ( .D(n2469), .CLK(clk), .RSTB(n3664), .Q(elem20[9]), 
        .QN(n791) );
  DFFARX1 \elem20_reg[8]  ( .D(n2468), .CLK(clk), .RSTB(n3664), .Q(elem20[8]), 
        .QN(n792) );
  DFFARX1 \elem20_reg[7]  ( .D(n2467), .CLK(clk), .RSTB(n3664), .Q(elem20[7]), 
        .QN(n793) );
  DFFARX1 \elem20_reg[6]  ( .D(n2466), .CLK(clk), .RSTB(n3664), .Q(elem20[6]), 
        .QN(n794) );
  DFFARX1 \elem20_reg[5]  ( .D(n2465), .CLK(clk), .RSTB(n3664), .Q(elem20[5]), 
        .QN(n795) );
  DFFARX1 \elem20_reg[4]  ( .D(n2464), .CLK(clk), .RSTB(n3664), .Q(elem20[4]), 
        .QN(n796) );
  DFFARX1 \elem20_reg[3]  ( .D(n2463), .CLK(clk), .RSTB(n3664), .Q(elem20[3]), 
        .QN(n797) );
  DFFARX1 \elem20_reg[2]  ( .D(n2462), .CLK(clk), .RSTB(n3664), .Q(elem20[2]), 
        .QN(n798) );
  DFFARX1 \elem20_reg[1]  ( .D(n2461), .CLK(clk), .RSTB(n3664), .Q(elem20[1]), 
        .QN(n799) );
  DFFARX1 \elem20_reg[0]  ( .D(n2460), .CLK(clk), .RSTB(n3664), .Q(elem20[0]), 
        .QN(n800) );
  DFFARX1 \elem21_reg[31]  ( .D(n2459), .CLK(clk), .RSTB(n3663), .Q(elem21[31]), .QN(n801) );
  DFFARX1 \elem21_reg[30]  ( .D(n2458), .CLK(clk), .RSTB(n3663), .Q(elem21[30]), .QN(n802) );
  DFFARX1 \elem21_reg[29]  ( .D(n2457), .CLK(clk), .RSTB(n3663), .Q(elem21[29]), .QN(n803) );
  DFFARX1 \elem21_reg[28]  ( .D(n2456), .CLK(clk), .RSTB(n3663), .Q(elem21[28]), .QN(n804) );
  DFFARX1 \elem21_reg[27]  ( .D(n2455), .CLK(clk), .RSTB(n3663), .Q(elem21[27]), .QN(n805) );
  DFFARX1 \elem21_reg[26]  ( .D(n2454), .CLK(clk), .RSTB(n3663), .Q(elem21[26]), .QN(n806) );
  DFFARX1 \elem21_reg[25]  ( .D(n2453), .CLK(clk), .RSTB(n3663), .Q(elem21[25]), .QN(n807) );
  DFFARX1 \elem21_reg[24]  ( .D(n2452), .CLK(clk), .RSTB(n3663), .Q(elem21[24]), .QN(n808) );
  DFFARX1 \elem21_reg[23]  ( .D(n2451), .CLK(clk), .RSTB(n3663), .Q(elem21[23]), .QN(n809) );
  DFFARX1 \elem21_reg[22]  ( .D(n2450), .CLK(clk), .RSTB(n3663), .Q(elem21[22]), .QN(n810) );
  DFFARX1 \elem21_reg[21]  ( .D(n2449), .CLK(clk), .RSTB(n3663), .Q(elem21[21]), .QN(n811) );
  DFFARX1 \elem21_reg[20]  ( .D(n2448), .CLK(clk), .RSTB(n3663), .Q(elem21[20]), .QN(n812) );
  DFFARX1 \elem21_reg[19]  ( .D(n2447), .CLK(clk), .RSTB(n3662), .Q(elem21[19]), .QN(n813) );
  DFFARX1 \elem21_reg[18]  ( .D(n2446), .CLK(clk), .RSTB(n3662), .Q(elem21[18]), .QN(n814) );
  DFFARX1 \elem21_reg[17]  ( .D(n2445), .CLK(clk), .RSTB(n3662), .Q(elem21[17]), .QN(n815) );
  DFFARX1 \elem21_reg[16]  ( .D(n2444), .CLK(clk), .RSTB(n3662), .Q(elem21[16]), .QN(n816) );
  DFFARX1 \elem21_reg[15]  ( .D(n2443), .CLK(clk), .RSTB(n3662), .Q(elem21[15]), .QN(n817) );
  DFFARX1 \elem21_reg[14]  ( .D(n2442), .CLK(clk), .RSTB(n3662), .Q(elem21[14]), .QN(n818) );
  DFFARX1 \elem21_reg[13]  ( .D(n2441), .CLK(clk), .RSTB(n3662), .Q(elem21[13]), .QN(n819) );
  DFFARX1 \elem21_reg[12]  ( .D(n2440), .CLK(clk), .RSTB(n3662), .Q(elem21[12]), .QN(n820) );
  DFFARX1 \elem21_reg[11]  ( .D(n2439), .CLK(clk), .RSTB(n3662), .Q(elem21[11]), .QN(n821) );
  DFFARX1 \elem21_reg[10]  ( .D(n2438), .CLK(clk), .RSTB(n3662), .Q(elem21[10]), .QN(n822) );
  DFFARX1 \elem21_reg[9]  ( .D(n2437), .CLK(clk), .RSTB(n3662), .Q(elem21[9]), 
        .QN(n823) );
  DFFARX1 \elem21_reg[8]  ( .D(n2436), .CLK(clk), .RSTB(n3662), .Q(elem21[8]), 
        .QN(n824) );
  DFFARX1 \elem21_reg[7]  ( .D(n2435), .CLK(clk), .RSTB(n3661), .Q(elem21[7]), 
        .QN(n825) );
  DFFARX1 \elem21_reg[6]  ( .D(n2434), .CLK(clk), .RSTB(n3661), .Q(elem21[6]), 
        .QN(n826) );
  DFFARX1 \elem21_reg[5]  ( .D(n2433), .CLK(clk), .RSTB(n3661), .Q(elem21[5]), 
        .QN(n827) );
  DFFARX1 \elem21_reg[4]  ( .D(n2432), .CLK(clk), .RSTB(n3661), .Q(elem21[4]), 
        .QN(n828) );
  DFFARX1 \elem21_reg[3]  ( .D(n2431), .CLK(clk), .RSTB(n3661), .Q(elem21[3]), 
        .QN(n829) );
  DFFARX1 \elem21_reg[2]  ( .D(n2430), .CLK(clk), .RSTB(n3661), .Q(elem21[2]), 
        .QN(n830) );
  DFFARX1 \elem21_reg[1]  ( .D(n2429), .CLK(clk), .RSTB(n3661), .Q(elem21[1]), 
        .QN(n831) );
  DFFARX1 \elem21_reg[0]  ( .D(n2428), .CLK(clk), .RSTB(n3661), .Q(elem21[0]), 
        .QN(n832) );
  DFFARX1 \elem22_reg[31]  ( .D(n2427), .CLK(clk), .RSTB(n3661), .Q(elem22[31]), .QN(n833) );
  DFFARX1 \elem22_reg[30]  ( .D(n2426), .CLK(clk), .RSTB(n3661), .Q(elem22[30]), .QN(n834) );
  DFFARX1 \elem22_reg[29]  ( .D(n2425), .CLK(clk), .RSTB(n3661), .Q(elem22[29]), .QN(n835) );
  DFFARX1 \elem22_reg[28]  ( .D(n2424), .CLK(clk), .RSTB(n3661), .Q(elem22[28]), .QN(n836) );
  DFFARX1 \elem22_reg[27]  ( .D(n2423), .CLK(clk), .RSTB(n3660), .Q(elem22[27]), .QN(n837) );
  DFFARX1 \elem22_reg[26]  ( .D(n2422), .CLK(clk), .RSTB(n3660), .Q(elem22[26]), .QN(n838) );
  DFFARX1 \elem22_reg[25]  ( .D(n2421), .CLK(clk), .RSTB(n3660), .Q(elem22[25]), .QN(n839) );
  DFFARX1 \elem22_reg[24]  ( .D(n2420), .CLK(clk), .RSTB(n3660), .Q(elem22[24]), .QN(n840) );
  DFFARX1 \elem22_reg[23]  ( .D(n2419), .CLK(clk), .RSTB(n3660), .Q(elem22[23]), .QN(n841) );
  DFFARX1 \elem22_reg[22]  ( .D(n2418), .CLK(clk), .RSTB(n3660), .Q(elem22[22]), .QN(n842) );
  DFFARX1 \elem22_reg[21]  ( .D(n2417), .CLK(clk), .RSTB(n3660), .Q(elem22[21]), .QN(n843) );
  DFFARX1 \elem22_reg[20]  ( .D(n2416), .CLK(clk), .RSTB(n3660), .Q(elem22[20]), .QN(n844) );
  DFFARX1 \elem22_reg[19]  ( .D(n2415), .CLK(clk), .RSTB(n3660), .Q(elem22[19]), .QN(n845) );
  DFFARX1 \elem22_reg[18]  ( .D(n2414), .CLK(clk), .RSTB(n3660), .Q(elem22[18]), .QN(n846) );
  DFFARX1 \elem22_reg[17]  ( .D(n2413), .CLK(clk), .RSTB(n3660), .Q(elem22[17]), .QN(n847) );
  DFFARX1 \elem22_reg[16]  ( .D(n2412), .CLK(clk), .RSTB(n3660), .Q(elem22[16]), .QN(n848) );
  DFFARX1 \elem22_reg[15]  ( .D(n2411), .CLK(clk), .RSTB(n3659), .Q(elem22[15]), .QN(n849) );
  DFFARX1 \elem22_reg[14]  ( .D(n2410), .CLK(clk), .RSTB(n3659), .Q(elem22[14]), .QN(n850) );
  DFFARX1 \elem22_reg[13]  ( .D(n2409), .CLK(clk), .RSTB(n3659), .Q(elem22[13]), .QN(n851) );
  DFFARX1 \elem22_reg[12]  ( .D(n2408), .CLK(clk), .RSTB(n3659), .Q(elem22[12]), .QN(n852) );
  DFFARX1 \elem22_reg[11]  ( .D(n2407), .CLK(clk), .RSTB(n3659), .Q(elem22[11]), .QN(n853) );
  DFFARX1 \elem22_reg[10]  ( .D(n2406), .CLK(clk), .RSTB(n3659), .Q(elem22[10]), .QN(n854) );
  DFFARX1 \elem22_reg[9]  ( .D(n2405), .CLK(clk), .RSTB(n3659), .Q(elem22[9]), 
        .QN(n855) );
  DFFARX1 \elem22_reg[8]  ( .D(n2404), .CLK(clk), .RSTB(n3659), .Q(elem22[8]), 
        .QN(n856) );
  DFFARX1 \elem22_reg[7]  ( .D(n2403), .CLK(clk), .RSTB(n3659), .Q(elem22[7]), 
        .QN(n857) );
  DFFARX1 \elem22_reg[6]  ( .D(n2402), .CLK(clk), .RSTB(n3659), .Q(elem22[6]), 
        .QN(n858) );
  DFFARX1 \elem22_reg[5]  ( .D(n2401), .CLK(clk), .RSTB(n3659), .Q(elem22[5]), 
        .QN(n859) );
  DFFARX1 \elem22_reg[4]  ( .D(n2400), .CLK(clk), .RSTB(n3659), .Q(elem22[4]), 
        .QN(n860) );
  DFFARX1 \elem22_reg[3]  ( .D(n2399), .CLK(clk), .RSTB(n3658), .Q(elem22[3]), 
        .QN(n861) );
  DFFARX1 \elem22_reg[2]  ( .D(n2398), .CLK(clk), .RSTB(n3658), .Q(elem22[2]), 
        .QN(n862) );
  DFFARX1 \elem22_reg[1]  ( .D(n2397), .CLK(clk), .RSTB(n3658), .Q(elem22[1]), 
        .QN(n863) );
  DFFARX1 \elem22_reg[0]  ( .D(n2396), .CLK(clk), .RSTB(n3658), .Q(elem22[0]), 
        .QN(n864) );
  DFFARX1 \elem23_reg[31]  ( .D(n2395), .CLK(clk), .RSTB(n3658), .Q(elem23[31]), .QN(n865) );
  DFFARX1 \elem23_reg[30]  ( .D(n2394), .CLK(clk), .RSTB(n3658), .Q(elem23[30]), .QN(n866) );
  DFFARX1 \elem23_reg[29]  ( .D(n2393), .CLK(clk), .RSTB(n3658), .Q(elem23[29]), .QN(n867) );
  DFFARX1 \elem23_reg[28]  ( .D(n2392), .CLK(clk), .RSTB(n3658), .Q(elem23[28]), .QN(n868) );
  DFFARX1 \elem23_reg[27]  ( .D(n2391), .CLK(clk), .RSTB(n3658), .Q(elem23[27]), .QN(n869) );
  DFFARX1 \elem23_reg[26]  ( .D(n2390), .CLK(clk), .RSTB(n3658), .Q(elem23[26]), .QN(n870) );
  DFFARX1 \elem23_reg[25]  ( .D(n2389), .CLK(clk), .RSTB(n3658), .Q(elem23[25]), .QN(n871) );
  DFFARX1 \elem23_reg[24]  ( .D(n2388), .CLK(clk), .RSTB(n3658), .Q(elem23[24]), .QN(n872) );
  DFFARX1 \elem23_reg[23]  ( .D(n2387), .CLK(clk), .RSTB(n3657), .Q(elem23[23]), .QN(n873) );
  DFFARX1 \elem23_reg[22]  ( .D(n2386), .CLK(clk), .RSTB(n3657), .Q(elem23[22]), .QN(n874) );
  DFFARX1 \elem23_reg[21]  ( .D(n2385), .CLK(clk), .RSTB(n3657), .Q(elem23[21]), .QN(n875) );
  DFFARX1 \elem23_reg[20]  ( .D(n2384), .CLK(clk), .RSTB(n3657), .Q(elem23[20]), .QN(n876) );
  DFFARX1 \elem23_reg[19]  ( .D(n2383), .CLK(clk), .RSTB(n3657), .Q(elem23[19]), .QN(n877) );
  DFFARX1 \elem23_reg[18]  ( .D(n2382), .CLK(clk), .RSTB(n3657), .Q(elem23[18]), .QN(n878) );
  DFFARX1 \elem23_reg[17]  ( .D(n2381), .CLK(clk), .RSTB(n3657), .Q(elem23[17]), .QN(n879) );
  DFFARX1 \elem23_reg[16]  ( .D(n2380), .CLK(clk), .RSTB(n3657), .Q(elem23[16]), .QN(n880) );
  DFFARX1 \elem23_reg[15]  ( .D(n2379), .CLK(clk), .RSTB(n3657), .Q(elem23[15]), .QN(n881) );
  DFFARX1 \elem23_reg[14]  ( .D(n2378), .CLK(clk), .RSTB(n3657), .Q(elem23[14]), .QN(n882) );
  DFFARX1 \elem23_reg[13]  ( .D(n2377), .CLK(clk), .RSTB(n3657), .Q(elem23[13]), .QN(n883) );
  DFFARX1 \elem23_reg[12]  ( .D(n2376), .CLK(clk), .RSTB(n3657), .Q(elem23[12]), .QN(n884) );
  DFFARX1 \elem23_reg[11]  ( .D(n2375), .CLK(clk), .RSTB(n3656), .Q(elem23[11]), .QN(n885) );
  DFFARX1 \elem23_reg[10]  ( .D(n2374), .CLK(clk), .RSTB(n3656), .Q(elem23[10]), .QN(n886) );
  DFFARX1 \elem23_reg[9]  ( .D(n2373), .CLK(clk), .RSTB(n3656), .Q(elem23[9]), 
        .QN(n887) );
  DFFARX1 \elem23_reg[8]  ( .D(n2372), .CLK(clk), .RSTB(n3656), .Q(elem23[8]), 
        .QN(n888) );
  DFFARX1 \elem23_reg[7]  ( .D(n2371), .CLK(clk), .RSTB(n3656), .Q(elem23[7]), 
        .QN(n889) );
  DFFARX1 \elem23_reg[6]  ( .D(n2370), .CLK(clk), .RSTB(n3656), .Q(elem23[6]), 
        .QN(n890) );
  DFFARX1 \elem23_reg[5]  ( .D(n2369), .CLK(clk), .RSTB(n3656), .Q(elem23[5]), 
        .QN(n891) );
  DFFARX1 \elem23_reg[4]  ( .D(n2368), .CLK(clk), .RSTB(n3656), .Q(elem23[4]), 
        .QN(n892) );
  DFFARX1 \elem23_reg[3]  ( .D(n2367), .CLK(clk), .RSTB(n3656), .Q(elem23[3]), 
        .QN(n893) );
  DFFARX1 \elem23_reg[2]  ( .D(n2366), .CLK(clk), .RSTB(n3656), .Q(elem23[2]), 
        .QN(n894) );
  DFFARX1 \elem23_reg[1]  ( .D(n2365), .CLK(clk), .RSTB(n3656), .Q(elem23[1]), 
        .QN(n895) );
  DFFARX1 \elem23_reg[0]  ( .D(n2364), .CLK(clk), .RSTB(n3656), .Q(elem23[0]), 
        .QN(n896) );
  DFFARX1 \elem24_reg[31]  ( .D(n2363), .CLK(clk), .RSTB(n3655), .Q(elem24[31]), .QN(n897) );
  DFFARX1 \elem24_reg[30]  ( .D(n2362), .CLK(clk), .RSTB(n3655), .Q(elem24[30]), .QN(n898) );
  DFFARX1 \elem24_reg[29]  ( .D(n2361), .CLK(clk), .RSTB(n3655), .Q(elem24[29]), .QN(n899) );
  DFFARX1 \elem24_reg[28]  ( .D(n2360), .CLK(clk), .RSTB(n3655), .Q(elem24[28]), .QN(n900) );
  DFFARX1 \elem24_reg[27]  ( .D(n2359), .CLK(clk), .RSTB(n3655), .Q(elem24[27]), .QN(n901) );
  DFFARX1 \elem24_reg[26]  ( .D(n2358), .CLK(clk), .RSTB(n3655), .Q(elem24[26]), .QN(n902) );
  DFFARX1 \elem24_reg[25]  ( .D(n2357), .CLK(clk), .RSTB(n3655), .Q(elem24[25]), .QN(n903) );
  DFFARX1 \elem24_reg[24]  ( .D(n2356), .CLK(clk), .RSTB(n3655), .Q(elem24[24]), .QN(n904) );
  DFFARX1 \elem24_reg[23]  ( .D(n2355), .CLK(clk), .RSTB(n3655), .Q(elem24[23]), .QN(n905) );
  DFFARX1 \elem24_reg[22]  ( .D(n2354), .CLK(clk), .RSTB(n3655), .Q(elem24[22]), .QN(n906) );
  DFFARX1 \elem24_reg[21]  ( .D(n2353), .CLK(clk), .RSTB(n3655), .Q(elem24[21]), .QN(n907) );
  DFFARX1 \elem24_reg[20]  ( .D(n2352), .CLK(clk), .RSTB(n3655), .Q(elem24[20]), .QN(n908) );
  DFFARX1 \elem24_reg[19]  ( .D(n2351), .CLK(clk), .RSTB(n3654), .Q(elem24[19]), .QN(n909) );
  DFFARX1 \elem24_reg[18]  ( .D(n2350), .CLK(clk), .RSTB(n3654), .Q(elem24[18]), .QN(n910) );
  DFFARX1 \elem24_reg[17]  ( .D(n2349), .CLK(clk), .RSTB(n3654), .Q(elem24[17]), .QN(n911) );
  DFFARX1 \elem24_reg[16]  ( .D(n2348), .CLK(clk), .RSTB(n3654), .Q(elem24[16]), .QN(n912) );
  DFFARX1 \elem24_reg[15]  ( .D(n2347), .CLK(clk), .RSTB(n3654), .Q(elem24[15]), .QN(n913) );
  DFFARX1 \elem24_reg[14]  ( .D(n2346), .CLK(clk), .RSTB(n3654), .Q(elem24[14]), .QN(n914) );
  DFFARX1 \elem24_reg[13]  ( .D(n2345), .CLK(clk), .RSTB(n3654), .Q(elem24[13]), .QN(n915) );
  DFFARX1 \elem24_reg[12]  ( .D(n2344), .CLK(clk), .RSTB(n3654), .Q(elem24[12]), .QN(n916) );
  DFFARX1 \elem24_reg[11]  ( .D(n2343), .CLK(clk), .RSTB(n3654), .Q(elem24[11]), .QN(n917) );
  DFFARX1 \elem24_reg[10]  ( .D(n2342), .CLK(clk), .RSTB(n3654), .Q(elem24[10]), .QN(n918) );
  DFFARX1 \elem24_reg[9]  ( .D(n2341), .CLK(clk), .RSTB(n3654), .Q(elem24[9]), 
        .QN(n919) );
  DFFARX1 \elem24_reg[8]  ( .D(n2340), .CLK(clk), .RSTB(n3654), .Q(elem24[8]), 
        .QN(n920) );
  DFFARX1 \elem24_reg[7]  ( .D(n2339), .CLK(clk), .RSTB(n3653), .Q(elem24[7]), 
        .QN(n921) );
  DFFARX1 \elem24_reg[6]  ( .D(n2338), .CLK(clk), .RSTB(n3653), .Q(elem24[6]), 
        .QN(n922) );
  DFFARX1 \elem24_reg[5]  ( .D(n2337), .CLK(clk), .RSTB(n3653), .Q(elem24[5]), 
        .QN(n923) );
  DFFARX1 \elem24_reg[4]  ( .D(n2336), .CLK(clk), .RSTB(n3653), .Q(elem24[4]), 
        .QN(n924) );
  DFFARX1 \elem24_reg[3]  ( .D(n2335), .CLK(clk), .RSTB(n3653), .Q(elem24[3]), 
        .QN(n925) );
  DFFARX1 \elem24_reg[2]  ( .D(n2334), .CLK(clk), .RSTB(n3653), .Q(elem24[2]), 
        .QN(n926) );
  DFFARX1 \elem24_reg[1]  ( .D(n2333), .CLK(clk), .RSTB(n3653), .Q(elem24[1]), 
        .QN(n927) );
  DFFARX1 \elem24_reg[0]  ( .D(n2332), .CLK(clk), .RSTB(n3653), .Q(elem24[0]), 
        .QN(n928) );
  DFFARX1 \elem25_reg[31]  ( .D(n2331), .CLK(clk), .RSTB(n3653), .Q(elem25[31]), .QN(n929) );
  DFFARX1 \elem25_reg[30]  ( .D(n2330), .CLK(clk), .RSTB(n3653), .Q(elem25[30]), .QN(n930) );
  DFFARX1 \elem25_reg[29]  ( .D(n2329), .CLK(clk), .RSTB(n3653), .Q(elem25[29]), .QN(n931) );
  DFFARX1 \elem25_reg[28]  ( .D(n2328), .CLK(clk), .RSTB(n3653), .Q(elem25[28]), .QN(n932) );
  DFFARX1 \elem25_reg[27]  ( .D(n2327), .CLK(clk), .RSTB(n3652), .Q(elem25[27]), .QN(n933) );
  DFFARX1 \elem25_reg[26]  ( .D(n2326), .CLK(clk), .RSTB(n3652), .Q(elem25[26]), .QN(n934) );
  DFFARX1 \elem25_reg[25]  ( .D(n2325), .CLK(clk), .RSTB(n3652), .Q(elem25[25]), .QN(n935) );
  DFFARX1 \elem25_reg[24]  ( .D(n2324), .CLK(clk), .RSTB(n3652), .Q(elem25[24]), .QN(n936) );
  DFFARX1 \elem25_reg[23]  ( .D(n2323), .CLK(clk), .RSTB(n3652), .Q(elem25[23]), .QN(n937) );
  DFFARX1 \elem25_reg[22]  ( .D(n2322), .CLK(clk), .RSTB(n3652), .Q(elem25[22]), .QN(n938) );
  DFFARX1 \elem25_reg[21]  ( .D(n2321), .CLK(clk), .RSTB(n3652), .Q(elem25[21]), .QN(n939) );
  DFFARX1 \elem25_reg[20]  ( .D(n2320), .CLK(clk), .RSTB(n3652), .Q(elem25[20]), .QN(n940) );
  DFFARX1 \elem25_reg[19]  ( .D(n2319), .CLK(clk), .RSTB(n3652), .Q(elem25[19]), .QN(n941) );
  DFFARX1 \elem25_reg[18]  ( .D(n2318), .CLK(clk), .RSTB(n3652), .Q(elem25[18]), .QN(n942) );
  DFFARX1 \elem25_reg[17]  ( .D(n2317), .CLK(clk), .RSTB(n3652), .Q(elem25[17]), .QN(n943) );
  DFFARX1 \elem25_reg[16]  ( .D(n2316), .CLK(clk), .RSTB(n3652), .Q(elem25[16]), .QN(n944) );
  DFFARX1 \elem25_reg[15]  ( .D(n2315), .CLK(clk), .RSTB(n3651), .Q(elem25[15]), .QN(n945) );
  DFFARX1 \elem25_reg[14]  ( .D(n2314), .CLK(clk), .RSTB(n3651), .Q(elem25[14]), .QN(n946) );
  DFFARX1 \elem25_reg[13]  ( .D(n2313), .CLK(clk), .RSTB(n3651), .Q(elem25[13]), .QN(n947) );
  DFFARX1 \elem25_reg[12]  ( .D(n2312), .CLK(clk), .RSTB(n3651), .Q(elem25[12]), .QN(n948) );
  DFFARX1 \elem25_reg[11]  ( .D(n2311), .CLK(clk), .RSTB(n3651), .Q(elem25[11]), .QN(n949) );
  DFFARX1 \elem25_reg[10]  ( .D(n2310), .CLK(clk), .RSTB(n3651), .Q(elem25[10]), .QN(n950) );
  DFFARX1 \elem25_reg[9]  ( .D(n2309), .CLK(clk), .RSTB(n3651), .Q(elem25[9]), 
        .QN(n951) );
  DFFARX1 \elem25_reg[8]  ( .D(n2308), .CLK(clk), .RSTB(n3651), .Q(elem25[8]), 
        .QN(n952) );
  DFFARX1 \elem25_reg[7]  ( .D(n2307), .CLK(clk), .RSTB(n3651), .Q(elem25[7]), 
        .QN(n953) );
  DFFARX1 \elem25_reg[6]  ( .D(n2306), .CLK(clk), .RSTB(n3651), .Q(elem25[6]), 
        .QN(n954) );
  DFFARX1 \elem25_reg[5]  ( .D(n2305), .CLK(clk), .RSTB(n3651), .Q(elem25[5]), 
        .QN(n955) );
  DFFARX1 \elem25_reg[4]  ( .D(n2304), .CLK(clk), .RSTB(n3651), .Q(elem25[4]), 
        .QN(n956) );
  DFFARX1 \elem25_reg[3]  ( .D(n2303), .CLK(clk), .RSTB(n3650), .Q(elem25[3]), 
        .QN(n957) );
  DFFARX1 \elem25_reg[2]  ( .D(n2302), .CLK(clk), .RSTB(n3650), .Q(elem25[2]), 
        .QN(n958) );
  DFFARX1 \elem25_reg[1]  ( .D(n2301), .CLK(clk), .RSTB(n3650), .Q(elem25[1]), 
        .QN(n959) );
  DFFARX1 \elem25_reg[0]  ( .D(n2300), .CLK(clk), .RSTB(n3650), .Q(elem25[0]), 
        .QN(n960) );
  DFFARX1 \elem26_reg[31]  ( .D(n2299), .CLK(clk), .RSTB(n3650), .Q(elem26[31]), .QN(n961) );
  DFFARX1 \elem26_reg[30]  ( .D(n2298), .CLK(clk), .RSTB(n3650), .Q(elem26[30]), .QN(n962) );
  DFFARX1 \elem26_reg[29]  ( .D(n2297), .CLK(clk), .RSTB(n3650), .Q(elem26[29]), .QN(n963) );
  DFFARX1 \elem26_reg[28]  ( .D(n2296), .CLK(clk), .RSTB(n3650), .Q(elem26[28]), .QN(n964) );
  DFFARX1 \elem26_reg[27]  ( .D(n2295), .CLK(clk), .RSTB(n3650), .Q(elem26[27]), .QN(n965) );
  DFFARX1 \elem26_reg[26]  ( .D(n2294), .CLK(clk), .RSTB(n3650), .Q(elem26[26]), .QN(n966) );
  DFFARX1 \elem26_reg[25]  ( .D(n2293), .CLK(clk), .RSTB(n3650), .Q(elem26[25]), .QN(n967) );
  DFFARX1 \elem26_reg[24]  ( .D(n2292), .CLK(clk), .RSTB(n3650), .Q(elem26[24]), .QN(n968) );
  DFFARX1 \elem26_reg[23]  ( .D(n2291), .CLK(clk), .RSTB(n3649), .Q(elem26[23]), .QN(n969) );
  DFFARX1 \elem26_reg[22]  ( .D(n2290), .CLK(clk), .RSTB(n3649), .Q(elem26[22]), .QN(n970) );
  DFFARX1 \elem26_reg[21]  ( .D(n2289), .CLK(clk), .RSTB(n3649), .Q(elem26[21]), .QN(n971) );
  DFFARX1 \elem26_reg[20]  ( .D(n2288), .CLK(clk), .RSTB(n3649), .Q(elem26[20]), .QN(n972) );
  DFFARX1 \elem26_reg[19]  ( .D(n2287), .CLK(clk), .RSTB(n3649), .Q(elem26[19]), .QN(n973) );
  DFFARX1 \elem26_reg[18]  ( .D(n2286), .CLK(clk), .RSTB(n3649), .Q(elem26[18]), .QN(n974) );
  DFFARX1 \elem26_reg[17]  ( .D(n2285), .CLK(clk), .RSTB(n3649), .Q(elem26[17]), .QN(n975) );
  DFFARX1 \elem26_reg[16]  ( .D(n2284), .CLK(clk), .RSTB(n3649), .Q(elem26[16]), .QN(n976) );
  DFFARX1 \elem26_reg[15]  ( .D(n2283), .CLK(clk), .RSTB(n3649), .Q(elem26[15]), .QN(n977) );
  DFFARX1 \elem26_reg[14]  ( .D(n2282), .CLK(clk), .RSTB(n3649), .Q(elem26[14]), .QN(n978) );
  DFFARX1 \elem26_reg[13]  ( .D(n2281), .CLK(clk), .RSTB(n3649), .Q(elem26[13]), .QN(n979) );
  DFFARX1 \elem26_reg[12]  ( .D(n2280), .CLK(clk), .RSTB(n3649), .Q(elem26[12]), .QN(n980) );
  DFFARX1 \elem26_reg[11]  ( .D(n2279), .CLK(clk), .RSTB(n3648), .Q(elem26[11]), .QN(n981) );
  DFFARX1 \elem26_reg[10]  ( .D(n2278), .CLK(clk), .RSTB(n3648), .Q(elem26[10]), .QN(n982) );
  DFFARX1 \elem26_reg[9]  ( .D(n2277), .CLK(clk), .RSTB(n3648), .Q(elem26[9]), 
        .QN(n983) );
  DFFARX1 \elem26_reg[8]  ( .D(n2276), .CLK(clk), .RSTB(n3648), .Q(elem26[8]), 
        .QN(n984) );
  DFFARX1 \elem26_reg[7]  ( .D(n2275), .CLK(clk), .RSTB(n3648), .Q(elem26[7]), 
        .QN(n985) );
  DFFARX1 \elem26_reg[6]  ( .D(n2274), .CLK(clk), .RSTB(n3648), .Q(elem26[6]), 
        .QN(n986) );
  DFFARX1 \elem26_reg[5]  ( .D(n2273), .CLK(clk), .RSTB(n3648), .Q(elem26[5]), 
        .QN(n987) );
  DFFARX1 \elem26_reg[4]  ( .D(n2272), .CLK(clk), .RSTB(n3648), .Q(elem26[4]), 
        .QN(n988) );
  DFFARX1 \elem26_reg[3]  ( .D(n2271), .CLK(clk), .RSTB(n3648), .Q(elem26[3]), 
        .QN(n989) );
  DFFARX1 \elem26_reg[2]  ( .D(n2270), .CLK(clk), .RSTB(n3648), .Q(elem26[2]), 
        .QN(n990) );
  DFFARX1 \elem26_reg[1]  ( .D(n2269), .CLK(clk), .RSTB(n3648), .Q(elem26[1]), 
        .QN(n991) );
  DFFARX1 \elem26_reg[0]  ( .D(n2268), .CLK(clk), .RSTB(n3648), .Q(elem26[0]), 
        .QN(n992) );
  OR2X1 U164 ( .IN1(n1039), .IN2(n1040), .Q(rd_dataB[9]) );
  NAND4X0 U165 ( .IN1(n1041), .IN2(n1042), .IN3(n1043), .IN4(n1044), .QN(n1040) );
  OA221X1 U166 ( .IN1(n3549), .IN2(n535), .IN3(n3546), .IN4(n567), .IN5(n1047), 
        .Q(n1044) );
  OA22X1 U167 ( .IN1(n3543), .IN2(n631), .IN3(n3540), .IN4(n599), .Q(n1047) );
  OA221X1 U168 ( .IN1(n3537), .IN2(n407), .IN3(n3534), .IN4(n439), .IN5(n1052), 
        .Q(n1043) );
  OA22X1 U169 ( .IN1(n3531), .IN2(n503), .IN3(n3528), .IN4(n471), .Q(n1052) );
  OA221X1 U170 ( .IN1(n3525), .IN2(n279), .IN3(n3522), .IN4(n311), .IN5(n1057), 
        .Q(n1042) );
  OA22X1 U171 ( .IN1(n3519), .IN2(n375), .IN3(n3516), .IN4(n343), .Q(n1057) );
  OA222X1 U172 ( .IN1(n3513), .IN2(n183), .IN3(n3510), .IN4(n247), .IN5(n3507), 
        .IN6(n215), .Q(n1041) );
  NAND4X0 U173 ( .IN1(n1063), .IN2(n1064), .IN3(n1065), .IN4(n1066), .QN(n1039) );
  OA221X1 U174 ( .IN1(n3504), .IN2(n119), .IN3(n3501), .IN4(n87), .IN5(n1069), 
        .Q(n1066) );
  OA22X1 U175 ( .IN1(n3498), .IN2(n151), .IN3(n3495), .IN4(n55), .Q(n1069) );
  OA221X1 U176 ( .IN1(n3492), .IN2(n919), .IN3(n3489), .IN4(n951), .IN5(n1074), 
        .Q(n1065) );
  OA22X1 U177 ( .IN1(n3486), .IN2(n23), .IN3(n3483), .IN4(n983), .Q(n1074) );
  OA221X1 U178 ( .IN1(n3480), .IN2(n791), .IN3(n3477), .IN4(n823), .IN5(n1079), 
        .Q(n1064) );
  OA22X1 U179 ( .IN1(n3474), .IN2(n887), .IN3(n3471), .IN4(n855), .Q(n1079) );
  OA221X1 U180 ( .IN1(n3468), .IN2(n727), .IN3(n3465), .IN4(n759), .IN5(n1084), 
        .Q(n1063) );
  OA22X1 U181 ( .IN1(n3462), .IN2(n695), .IN3(n3459), .IN4(n663), .Q(n1084) );
  OR2X1 U182 ( .IN1(n1087), .IN2(n1088), .Q(rd_dataB[8]) );
  NAND4X0 U183 ( .IN1(n1089), .IN2(n1090), .IN3(n1091), .IN4(n1092), .QN(n1088) );
  OA221X1 U184 ( .IN1(n3549), .IN2(n536), .IN3(n3546), .IN4(n568), .IN5(n1093), 
        .Q(n1092) );
  OA22X1 U185 ( .IN1(n3543), .IN2(n632), .IN3(n3540), .IN4(n600), .Q(n1093) );
  OA221X1 U186 ( .IN1(n3537), .IN2(n408), .IN3(n3534), .IN4(n440), .IN5(n1094), 
        .Q(n1091) );
  OA22X1 U187 ( .IN1(n3531), .IN2(n504), .IN3(n3528), .IN4(n472), .Q(n1094) );
  OA221X1 U188 ( .IN1(n3525), .IN2(n280), .IN3(n3522), .IN4(n312), .IN5(n1095), 
        .Q(n1090) );
  OA22X1 U189 ( .IN1(n3519), .IN2(n376), .IN3(n3516), .IN4(n344), .Q(n1095) );
  OA222X1 U190 ( .IN1(n3513), .IN2(n184), .IN3(n3510), .IN4(n248), .IN5(n3507), 
        .IN6(n216), .Q(n1089) );
  NAND4X0 U191 ( .IN1(n1096), .IN2(n1097), .IN3(n1098), .IN4(n1099), .QN(n1087) );
  OA221X1 U192 ( .IN1(n3504), .IN2(n120), .IN3(n3501), .IN4(n88), .IN5(n1100), 
        .Q(n1099) );
  OA22X1 U193 ( .IN1(n3498), .IN2(n152), .IN3(n3495), .IN4(n56), .Q(n1100) );
  OA221X1 U194 ( .IN1(n3492), .IN2(n920), .IN3(n3489), .IN4(n952), .IN5(n1101), 
        .Q(n1098) );
  OA22X1 U195 ( .IN1(n3486), .IN2(n24), .IN3(n3483), .IN4(n984), .Q(n1101) );
  OA221X1 U196 ( .IN1(n3480), .IN2(n792), .IN3(n3477), .IN4(n824), .IN5(n1102), 
        .Q(n1097) );
  OA22X1 U197 ( .IN1(n3474), .IN2(n888), .IN3(n3471), .IN4(n856), .Q(n1102) );
  OA221X1 U198 ( .IN1(n3468), .IN2(n728), .IN3(n3465), .IN4(n760), .IN5(n1103), 
        .Q(n1096) );
  OA22X1 U199 ( .IN1(n3462), .IN2(n696), .IN3(n3459), .IN4(n664), .Q(n1103) );
  OR2X1 U200 ( .IN1(n1104), .IN2(n1105), .Q(rd_dataB[7]) );
  NAND4X0 U201 ( .IN1(n1106), .IN2(n1107), .IN3(n1108), .IN4(n1109), .QN(n1105) );
  OA221X1 U202 ( .IN1(n3549), .IN2(n537), .IN3(n3546), .IN4(n569), .IN5(n1110), 
        .Q(n1109) );
  OA22X1 U203 ( .IN1(n3543), .IN2(n633), .IN3(n3540), .IN4(n601), .Q(n1110) );
  OA221X1 U204 ( .IN1(n3537), .IN2(n409), .IN3(n3534), .IN4(n441), .IN5(n1111), 
        .Q(n1108) );
  OA22X1 U205 ( .IN1(n3531), .IN2(n505), .IN3(n3528), .IN4(n473), .Q(n1111) );
  OA221X1 U206 ( .IN1(n3525), .IN2(n281), .IN3(n3522), .IN4(n313), .IN5(n1112), 
        .Q(n1107) );
  OA22X1 U207 ( .IN1(n3519), .IN2(n377), .IN3(n3516), .IN4(n345), .Q(n1112) );
  OA222X1 U208 ( .IN1(n3513), .IN2(n185), .IN3(n3510), .IN4(n249), .IN5(n3507), 
        .IN6(n217), .Q(n1106) );
  NAND4X0 U209 ( .IN1(n1113), .IN2(n1114), .IN3(n1115), .IN4(n1116), .QN(n1104) );
  OA221X1 U210 ( .IN1(n3504), .IN2(n121), .IN3(n3501), .IN4(n89), .IN5(n1117), 
        .Q(n1116) );
  OA22X1 U211 ( .IN1(n3498), .IN2(n153), .IN3(n3495), .IN4(n57), .Q(n1117) );
  OA221X1 U212 ( .IN1(n3492), .IN2(n921), .IN3(n3489), .IN4(n953), .IN5(n1118), 
        .Q(n1115) );
  OA22X1 U213 ( .IN1(n3486), .IN2(n25), .IN3(n3483), .IN4(n985), .Q(n1118) );
  OA221X1 U214 ( .IN1(n3480), .IN2(n793), .IN3(n3477), .IN4(n825), .IN5(n1119), 
        .Q(n1114) );
  OA22X1 U215 ( .IN1(n3474), .IN2(n889), .IN3(n3471), .IN4(n857), .Q(n1119) );
  OA221X1 U216 ( .IN1(n3468), .IN2(n729), .IN3(n3465), .IN4(n761), .IN5(n1120), 
        .Q(n1113) );
  OA22X1 U217 ( .IN1(n3462), .IN2(n697), .IN3(n3459), .IN4(n665), .Q(n1120) );
  OR2X1 U218 ( .IN1(n1121), .IN2(n1122), .Q(rd_dataB[6]) );
  NAND4X0 U219 ( .IN1(n1123), .IN2(n1124), .IN3(n1125), .IN4(n1126), .QN(n1122) );
  OA221X1 U220 ( .IN1(n3549), .IN2(n538), .IN3(n3546), .IN4(n570), .IN5(n1127), 
        .Q(n1126) );
  OA22X1 U221 ( .IN1(n3543), .IN2(n634), .IN3(n3540), .IN4(n602), .Q(n1127) );
  OA221X1 U222 ( .IN1(n3537), .IN2(n410), .IN3(n3534), .IN4(n442), .IN5(n1128), 
        .Q(n1125) );
  OA22X1 U223 ( .IN1(n3531), .IN2(n506), .IN3(n3528), .IN4(n474), .Q(n1128) );
  OA221X1 U224 ( .IN1(n3525), .IN2(n282), .IN3(n3522), .IN4(n314), .IN5(n1129), 
        .Q(n1124) );
  OA22X1 U225 ( .IN1(n3519), .IN2(n378), .IN3(n3516), .IN4(n346), .Q(n1129) );
  OA222X1 U226 ( .IN1(n3513), .IN2(n186), .IN3(n3510), .IN4(n250), .IN5(n3507), 
        .IN6(n218), .Q(n1123) );
  NAND4X0 U227 ( .IN1(n1130), .IN2(n1131), .IN3(n1132), .IN4(n1133), .QN(n1121) );
  OA221X1 U228 ( .IN1(n3504), .IN2(n122), .IN3(n3501), .IN4(n90), .IN5(n1134), 
        .Q(n1133) );
  OA22X1 U229 ( .IN1(n3498), .IN2(n154), .IN3(n3495), .IN4(n58), .Q(n1134) );
  OA221X1 U230 ( .IN1(n3492), .IN2(n922), .IN3(n3489), .IN4(n954), .IN5(n1135), 
        .Q(n1132) );
  OA22X1 U231 ( .IN1(n3486), .IN2(n26), .IN3(n3483), .IN4(n986), .Q(n1135) );
  OA221X1 U232 ( .IN1(n3480), .IN2(n794), .IN3(n3477), .IN4(n826), .IN5(n1136), 
        .Q(n1131) );
  OA22X1 U233 ( .IN1(n3474), .IN2(n890), .IN3(n3471), .IN4(n858), .Q(n1136) );
  OA221X1 U234 ( .IN1(n3468), .IN2(n730), .IN3(n3465), .IN4(n762), .IN5(n1137), 
        .Q(n1130) );
  OA22X1 U235 ( .IN1(n3462), .IN2(n698), .IN3(n3459), .IN4(n666), .Q(n1137) );
  OR2X1 U236 ( .IN1(n1138), .IN2(n1139), .Q(rd_dataB[5]) );
  NAND4X0 U237 ( .IN1(n1140), .IN2(n1141), .IN3(n1142), .IN4(n1143), .QN(n1139) );
  OA221X1 U238 ( .IN1(n3549), .IN2(n539), .IN3(n3546), .IN4(n571), .IN5(n1144), 
        .Q(n1143) );
  OA22X1 U239 ( .IN1(n3543), .IN2(n635), .IN3(n3540), .IN4(n603), .Q(n1144) );
  OA221X1 U240 ( .IN1(n3537), .IN2(n411), .IN3(n3534), .IN4(n443), .IN5(n1145), 
        .Q(n1142) );
  OA22X1 U241 ( .IN1(n3531), .IN2(n507), .IN3(n3528), .IN4(n475), .Q(n1145) );
  OA221X1 U242 ( .IN1(n3525), .IN2(n283), .IN3(n3522), .IN4(n315), .IN5(n1146), 
        .Q(n1141) );
  OA22X1 U243 ( .IN1(n3519), .IN2(n379), .IN3(n3516), .IN4(n347), .Q(n1146) );
  OA222X1 U244 ( .IN1(n3513), .IN2(n187), .IN3(n3510), .IN4(n251), .IN5(n3507), 
        .IN6(n219), .Q(n1140) );
  NAND4X0 U245 ( .IN1(n1147), .IN2(n1148), .IN3(n1149), .IN4(n1150), .QN(n1138) );
  OA221X1 U246 ( .IN1(n3504), .IN2(n123), .IN3(n3501), .IN4(n91), .IN5(n1151), 
        .Q(n1150) );
  OA22X1 U247 ( .IN1(n3498), .IN2(n155), .IN3(n3495), .IN4(n59), .Q(n1151) );
  OA221X1 U248 ( .IN1(n3492), .IN2(n923), .IN3(n3489), .IN4(n955), .IN5(n1152), 
        .Q(n1149) );
  OA22X1 U249 ( .IN1(n3486), .IN2(n27), .IN3(n3483), .IN4(n987), .Q(n1152) );
  OA221X1 U250 ( .IN1(n3480), .IN2(n795), .IN3(n3477), .IN4(n827), .IN5(n1153), 
        .Q(n1148) );
  OA22X1 U251 ( .IN1(n3474), .IN2(n891), .IN3(n3471), .IN4(n859), .Q(n1153) );
  OA221X1 U252 ( .IN1(n3468), .IN2(n731), .IN3(n3465), .IN4(n763), .IN5(n1154), 
        .Q(n1147) );
  OA22X1 U253 ( .IN1(n3462), .IN2(n699), .IN3(n3459), .IN4(n667), .Q(n1154) );
  OR2X1 U254 ( .IN1(n1155), .IN2(n1156), .Q(rd_dataB[4]) );
  NAND4X0 U255 ( .IN1(n1157), .IN2(n1158), .IN3(n1159), .IN4(n1160), .QN(n1156) );
  OA221X1 U256 ( .IN1(n3549), .IN2(n540), .IN3(n3546), .IN4(n572), .IN5(n1161), 
        .Q(n1160) );
  OA22X1 U257 ( .IN1(n3543), .IN2(n636), .IN3(n3540), .IN4(n604), .Q(n1161) );
  OA221X1 U258 ( .IN1(n3537), .IN2(n412), .IN3(n3534), .IN4(n444), .IN5(n1162), 
        .Q(n1159) );
  OA22X1 U259 ( .IN1(n3531), .IN2(n508), .IN3(n3528), .IN4(n476), .Q(n1162) );
  OA221X1 U260 ( .IN1(n3525), .IN2(n284), .IN3(n3522), .IN4(n316), .IN5(n1163), 
        .Q(n1158) );
  OA22X1 U261 ( .IN1(n3519), .IN2(n380), .IN3(n3516), .IN4(n348), .Q(n1163) );
  OA222X1 U262 ( .IN1(n3513), .IN2(n188), .IN3(n3510), .IN4(n252), .IN5(n3507), 
        .IN6(n220), .Q(n1157) );
  NAND4X0 U263 ( .IN1(n1164), .IN2(n1165), .IN3(n1166), .IN4(n1167), .QN(n1155) );
  OA221X1 U264 ( .IN1(n3504), .IN2(n124), .IN3(n3501), .IN4(n92), .IN5(n1168), 
        .Q(n1167) );
  OA22X1 U265 ( .IN1(n3498), .IN2(n156), .IN3(n3495), .IN4(n60), .Q(n1168) );
  OA221X1 U266 ( .IN1(n3492), .IN2(n924), .IN3(n3489), .IN4(n956), .IN5(n1169), 
        .Q(n1166) );
  OA22X1 U267 ( .IN1(n3486), .IN2(n28), .IN3(n3483), .IN4(n988), .Q(n1169) );
  OA221X1 U268 ( .IN1(n3480), .IN2(n796), .IN3(n3477), .IN4(n828), .IN5(n1170), 
        .Q(n1165) );
  OA22X1 U269 ( .IN1(n3474), .IN2(n892), .IN3(n3471), .IN4(n860), .Q(n1170) );
  OA221X1 U270 ( .IN1(n3468), .IN2(n732), .IN3(n3465), .IN4(n764), .IN5(n1171), 
        .Q(n1164) );
  OA22X1 U271 ( .IN1(n3462), .IN2(n700), .IN3(n3459), .IN4(n668), .Q(n1171) );
  OR2X1 U272 ( .IN1(n1172), .IN2(n1173), .Q(rd_dataB[3]) );
  NAND4X0 U273 ( .IN1(n1174), .IN2(n1175), .IN3(n1176), .IN4(n1177), .QN(n1173) );
  OA221X1 U274 ( .IN1(n3549), .IN2(n541), .IN3(n3546), .IN4(n573), .IN5(n1178), 
        .Q(n1177) );
  OA22X1 U275 ( .IN1(n3543), .IN2(n637), .IN3(n3540), .IN4(n605), .Q(n1178) );
  OA221X1 U276 ( .IN1(n3537), .IN2(n413), .IN3(n3534), .IN4(n445), .IN5(n1179), 
        .Q(n1176) );
  OA22X1 U277 ( .IN1(n3531), .IN2(n509), .IN3(n3528), .IN4(n477), .Q(n1179) );
  OA221X1 U278 ( .IN1(n3525), .IN2(n285), .IN3(n3522), .IN4(n317), .IN5(n1180), 
        .Q(n1175) );
  OA22X1 U279 ( .IN1(n3519), .IN2(n381), .IN3(n3516), .IN4(n349), .Q(n1180) );
  OA222X1 U280 ( .IN1(n3513), .IN2(n189), .IN3(n3510), .IN4(n253), .IN5(n3507), 
        .IN6(n221), .Q(n1174) );
  NAND4X0 U281 ( .IN1(n1181), .IN2(n1182), .IN3(n1183), .IN4(n1184), .QN(n1172) );
  OA221X1 U282 ( .IN1(n3504), .IN2(n125), .IN3(n3501), .IN4(n93), .IN5(n1185), 
        .Q(n1184) );
  OA22X1 U283 ( .IN1(n3498), .IN2(n157), .IN3(n3495), .IN4(n61), .Q(n1185) );
  OA221X1 U284 ( .IN1(n3492), .IN2(n925), .IN3(n3489), .IN4(n957), .IN5(n1186), 
        .Q(n1183) );
  OA22X1 U285 ( .IN1(n3486), .IN2(n29), .IN3(n3483), .IN4(n989), .Q(n1186) );
  OA221X1 U286 ( .IN1(n3480), .IN2(n797), .IN3(n3477), .IN4(n829), .IN5(n1187), 
        .Q(n1182) );
  OA22X1 U287 ( .IN1(n3474), .IN2(n893), .IN3(n3471), .IN4(n861), .Q(n1187) );
  OA221X1 U288 ( .IN1(n3468), .IN2(n733), .IN3(n3465), .IN4(n765), .IN5(n1188), 
        .Q(n1181) );
  OA22X1 U289 ( .IN1(n3462), .IN2(n701), .IN3(n3459), .IN4(n669), .Q(n1188) );
  OR2X1 U290 ( .IN1(n1189), .IN2(n1190), .Q(rd_dataB[31]) );
  NAND4X0 U291 ( .IN1(n1191), .IN2(n1192), .IN3(n1193), .IN4(n1194), .QN(n1190) );
  OA221X1 U292 ( .IN1(n3549), .IN2(n513), .IN3(n3546), .IN4(n545), .IN5(n1195), 
        .Q(n1194) );
  OA22X1 U293 ( .IN1(n3543), .IN2(n609), .IN3(n3540), .IN4(n577), .Q(n1195) );
  OA221X1 U294 ( .IN1(n3537), .IN2(n385), .IN3(n3534), .IN4(n417), .IN5(n1196), 
        .Q(n1193) );
  OA22X1 U295 ( .IN1(n3531), .IN2(n481), .IN3(n3528), .IN4(n449), .Q(n1196) );
  OA221X1 U296 ( .IN1(n3525), .IN2(n257), .IN3(n3522), .IN4(n289), .IN5(n1197), 
        .Q(n1192) );
  OA22X1 U297 ( .IN1(n3519), .IN2(n353), .IN3(n3516), .IN4(n321), .Q(n1197) );
  OA222X1 U298 ( .IN1(n3513), .IN2(n161), .IN3(n3510), .IN4(n225), .IN5(n3507), 
        .IN6(n193), .Q(n1191) );
  NAND4X0 U299 ( .IN1(n1198), .IN2(n1199), .IN3(n1200), .IN4(n1201), .QN(n1189) );
  OA221X1 U300 ( .IN1(n3504), .IN2(n97), .IN3(n3501), .IN4(n65), .IN5(n1202), 
        .Q(n1201) );
  OA22X1 U301 ( .IN1(n3498), .IN2(n129), .IN3(n3495), .IN4(n33), .Q(n1202) );
  OA221X1 U302 ( .IN1(n3492), .IN2(n897), .IN3(n3489), .IN4(n929), .IN5(n1203), 
        .Q(n1200) );
  OA22X1 U303 ( .IN1(n3486), .IN2(n1), .IN3(n3483), .IN4(n961), .Q(n1203) );
  OA221X1 U304 ( .IN1(n3480), .IN2(n769), .IN3(n3477), .IN4(n801), .IN5(n1204), 
        .Q(n1199) );
  OA22X1 U305 ( .IN1(n3474), .IN2(n865), .IN3(n3471), .IN4(n833), .Q(n1204) );
  OA221X1 U306 ( .IN1(n3468), .IN2(n705), .IN3(n3465), .IN4(n737), .IN5(n1205), 
        .Q(n1198) );
  OA22X1 U307 ( .IN1(n3462), .IN2(n673), .IN3(n3459), .IN4(n641), .Q(n1205) );
  OR2X1 U308 ( .IN1(n1206), .IN2(n1207), .Q(rd_dataB[30]) );
  NAND4X0 U309 ( .IN1(n1208), .IN2(n1209), .IN3(n1210), .IN4(n1211), .QN(n1207) );
  OA221X1 U310 ( .IN1(n3549), .IN2(n514), .IN3(n3546), .IN4(n546), .IN5(n1212), 
        .Q(n1211) );
  OA22X1 U311 ( .IN1(n3543), .IN2(n610), .IN3(n3540), .IN4(n578), .Q(n1212) );
  OA221X1 U312 ( .IN1(n3537), .IN2(n386), .IN3(n3534), .IN4(n418), .IN5(n1213), 
        .Q(n1210) );
  OA22X1 U313 ( .IN1(n3531), .IN2(n482), .IN3(n3528), .IN4(n450), .Q(n1213) );
  OA221X1 U314 ( .IN1(n3525), .IN2(n258), .IN3(n3522), .IN4(n290), .IN5(n1214), 
        .Q(n1209) );
  OA22X1 U315 ( .IN1(n3519), .IN2(n354), .IN3(n3516), .IN4(n322), .Q(n1214) );
  OA222X1 U316 ( .IN1(n3513), .IN2(n162), .IN3(n3510), .IN4(n226), .IN5(n3507), 
        .IN6(n194), .Q(n1208) );
  NAND4X0 U317 ( .IN1(n1215), .IN2(n1216), .IN3(n1217), .IN4(n1218), .QN(n1206) );
  OA221X1 U318 ( .IN1(n3504), .IN2(n98), .IN3(n3501), .IN4(n66), .IN5(n1219), 
        .Q(n1218) );
  OA22X1 U319 ( .IN1(n3498), .IN2(n130), .IN3(n3495), .IN4(n34), .Q(n1219) );
  OA221X1 U320 ( .IN1(n3492), .IN2(n898), .IN3(n3489), .IN4(n930), .IN5(n1220), 
        .Q(n1217) );
  OA22X1 U321 ( .IN1(n3486), .IN2(n2), .IN3(n3483), .IN4(n962), .Q(n1220) );
  OA221X1 U322 ( .IN1(n3480), .IN2(n770), .IN3(n3477), .IN4(n802), .IN5(n1221), 
        .Q(n1216) );
  OA22X1 U323 ( .IN1(n3474), .IN2(n866), .IN3(n3471), .IN4(n834), .Q(n1221) );
  OA221X1 U324 ( .IN1(n3468), .IN2(n706), .IN3(n3465), .IN4(n738), .IN5(n1222), 
        .Q(n1215) );
  OA22X1 U325 ( .IN1(n3462), .IN2(n674), .IN3(n3459), .IN4(n642), .Q(n1222) );
  OR2X1 U326 ( .IN1(n1223), .IN2(n1224), .Q(rd_dataB[2]) );
  NAND4X0 U327 ( .IN1(n1225), .IN2(n1226), .IN3(n1227), .IN4(n1228), .QN(n1224) );
  OA221X1 U328 ( .IN1(n3549), .IN2(n542), .IN3(n3546), .IN4(n574), .IN5(n1229), 
        .Q(n1228) );
  OA22X1 U329 ( .IN1(n3543), .IN2(n638), .IN3(n3540), .IN4(n606), .Q(n1229) );
  OA221X1 U330 ( .IN1(n3537), .IN2(n414), .IN3(n3534), .IN4(n446), .IN5(n1230), 
        .Q(n1227) );
  OA22X1 U331 ( .IN1(n3531), .IN2(n510), .IN3(n3528), .IN4(n478), .Q(n1230) );
  OA221X1 U332 ( .IN1(n3525), .IN2(n286), .IN3(n3522), .IN4(n318), .IN5(n1231), 
        .Q(n1226) );
  OA22X1 U333 ( .IN1(n3519), .IN2(n382), .IN3(n3516), .IN4(n350), .Q(n1231) );
  OA222X1 U334 ( .IN1(n3513), .IN2(n190), .IN3(n3510), .IN4(n254), .IN5(n3507), 
        .IN6(n222), .Q(n1225) );
  NAND4X0 U335 ( .IN1(n1232), .IN2(n1233), .IN3(n1234), .IN4(n1235), .QN(n1223) );
  OA221X1 U336 ( .IN1(n3504), .IN2(n126), .IN3(n3501), .IN4(n94), .IN5(n1236), 
        .Q(n1235) );
  OA22X1 U337 ( .IN1(n3498), .IN2(n158), .IN3(n3495), .IN4(n62), .Q(n1236) );
  OA221X1 U338 ( .IN1(n3492), .IN2(n926), .IN3(n3489), .IN4(n958), .IN5(n1237), 
        .Q(n1234) );
  OA22X1 U339 ( .IN1(n3486), .IN2(n30), .IN3(n3483), .IN4(n990), .Q(n1237) );
  OA221X1 U340 ( .IN1(n3480), .IN2(n798), .IN3(n3477), .IN4(n830), .IN5(n1238), 
        .Q(n1233) );
  OA22X1 U341 ( .IN1(n3474), .IN2(n894), .IN3(n3471), .IN4(n862), .Q(n1238) );
  OA221X1 U342 ( .IN1(n3468), .IN2(n734), .IN3(n3465), .IN4(n766), .IN5(n1239), 
        .Q(n1232) );
  OA22X1 U343 ( .IN1(n3462), .IN2(n702), .IN3(n3459), .IN4(n670), .Q(n1239) );
  OR2X1 U344 ( .IN1(n1240), .IN2(n1241), .Q(rd_dataB[29]) );
  NAND4X0 U345 ( .IN1(n1242), .IN2(n1243), .IN3(n1244), .IN4(n1245), .QN(n1241) );
  OA221X1 U346 ( .IN1(n3549), .IN2(n515), .IN3(n3546), .IN4(n547), .IN5(n1246), 
        .Q(n1245) );
  OA22X1 U347 ( .IN1(n3543), .IN2(n611), .IN3(n3540), .IN4(n579), .Q(n1246) );
  OA221X1 U348 ( .IN1(n3537), .IN2(n387), .IN3(n3534), .IN4(n419), .IN5(n1247), 
        .Q(n1244) );
  OA22X1 U349 ( .IN1(n3531), .IN2(n483), .IN3(n3528), .IN4(n451), .Q(n1247) );
  OA221X1 U350 ( .IN1(n3525), .IN2(n259), .IN3(n3522), .IN4(n291), .IN5(n1248), 
        .Q(n1243) );
  OA22X1 U351 ( .IN1(n3519), .IN2(n355), .IN3(n3516), .IN4(n323), .Q(n1248) );
  OA222X1 U352 ( .IN1(n3513), .IN2(n163), .IN3(n3510), .IN4(n227), .IN5(n3507), 
        .IN6(n195), .Q(n1242) );
  NAND4X0 U353 ( .IN1(n1249), .IN2(n1250), .IN3(n1251), .IN4(n1252), .QN(n1240) );
  OA221X1 U354 ( .IN1(n3504), .IN2(n99), .IN3(n3501), .IN4(n67), .IN5(n1253), 
        .Q(n1252) );
  OA22X1 U355 ( .IN1(n3498), .IN2(n131), .IN3(n3495), .IN4(n35), .Q(n1253) );
  OA221X1 U356 ( .IN1(n3492), .IN2(n899), .IN3(n3489), .IN4(n931), .IN5(n1254), 
        .Q(n1251) );
  OA22X1 U357 ( .IN1(n3486), .IN2(n3), .IN3(n3483), .IN4(n963), .Q(n1254) );
  OA221X1 U358 ( .IN1(n3480), .IN2(n771), .IN3(n3477), .IN4(n803), .IN5(n1255), 
        .Q(n1250) );
  OA22X1 U359 ( .IN1(n3474), .IN2(n867), .IN3(n3471), .IN4(n835), .Q(n1255) );
  OA221X1 U360 ( .IN1(n3468), .IN2(n707), .IN3(n3465), .IN4(n739), .IN5(n1256), 
        .Q(n1249) );
  OA22X1 U361 ( .IN1(n3462), .IN2(n675), .IN3(n3459), .IN4(n643), .Q(n1256) );
  OR2X1 U362 ( .IN1(n1257), .IN2(n1258), .Q(rd_dataB[28]) );
  NAND4X0 U363 ( .IN1(n1259), .IN2(n1260), .IN3(n1261), .IN4(n1262), .QN(n1258) );
  OA221X1 U364 ( .IN1(n3549), .IN2(n516), .IN3(n3546), .IN4(n548), .IN5(n1263), 
        .Q(n1262) );
  OA22X1 U365 ( .IN1(n3543), .IN2(n612), .IN3(n3540), .IN4(n580), .Q(n1263) );
  OA221X1 U366 ( .IN1(n3537), .IN2(n388), .IN3(n3534), .IN4(n420), .IN5(n1264), 
        .Q(n1261) );
  OA22X1 U367 ( .IN1(n3531), .IN2(n484), .IN3(n3528), .IN4(n452), .Q(n1264) );
  OA221X1 U368 ( .IN1(n3525), .IN2(n260), .IN3(n3522), .IN4(n292), .IN5(n1265), 
        .Q(n1260) );
  OA22X1 U369 ( .IN1(n3519), .IN2(n356), .IN3(n3516), .IN4(n324), .Q(n1265) );
  OA222X1 U370 ( .IN1(n3513), .IN2(n164), .IN3(n3510), .IN4(n228), .IN5(n3507), 
        .IN6(n196), .Q(n1259) );
  NAND4X0 U371 ( .IN1(n1266), .IN2(n1267), .IN3(n1268), .IN4(n1269), .QN(n1257) );
  OA221X1 U372 ( .IN1(n3504), .IN2(n100), .IN3(n3501), .IN4(n68), .IN5(n1270), 
        .Q(n1269) );
  OA22X1 U373 ( .IN1(n3498), .IN2(n132), .IN3(n3495), .IN4(n36), .Q(n1270) );
  OA221X1 U374 ( .IN1(n3492), .IN2(n900), .IN3(n3489), .IN4(n932), .IN5(n1271), 
        .Q(n1268) );
  OA22X1 U375 ( .IN1(n3486), .IN2(n4), .IN3(n3483), .IN4(n964), .Q(n1271) );
  OA221X1 U376 ( .IN1(n3480), .IN2(n772), .IN3(n3477), .IN4(n804), .IN5(n1272), 
        .Q(n1267) );
  OA22X1 U377 ( .IN1(n3474), .IN2(n868), .IN3(n3471), .IN4(n836), .Q(n1272) );
  OA221X1 U378 ( .IN1(n3468), .IN2(n708), .IN3(n3465), .IN4(n740), .IN5(n1273), 
        .Q(n1266) );
  OA22X1 U379 ( .IN1(n3462), .IN2(n676), .IN3(n3459), .IN4(n644), .Q(n1273) );
  OR2X1 U380 ( .IN1(n1274), .IN2(n1275), .Q(rd_dataB[27]) );
  NAND4X0 U381 ( .IN1(n1276), .IN2(n1277), .IN3(n1278), .IN4(n1279), .QN(n1275) );
  OA221X1 U382 ( .IN1(n3550), .IN2(n517), .IN3(n3547), .IN4(n549), .IN5(n1280), 
        .Q(n1279) );
  OA22X1 U383 ( .IN1(n3544), .IN2(n613), .IN3(n3541), .IN4(n581), .Q(n1280) );
  OA221X1 U384 ( .IN1(n3538), .IN2(n389), .IN3(n3535), .IN4(n421), .IN5(n1281), 
        .Q(n1278) );
  OA22X1 U385 ( .IN1(n3532), .IN2(n485), .IN3(n3529), .IN4(n453), .Q(n1281) );
  OA221X1 U386 ( .IN1(n3526), .IN2(n261), .IN3(n3523), .IN4(n293), .IN5(n1282), 
        .Q(n1277) );
  OA22X1 U387 ( .IN1(n3520), .IN2(n357), .IN3(n3517), .IN4(n325), .Q(n1282) );
  OA222X1 U388 ( .IN1(n3514), .IN2(n165), .IN3(n3511), .IN4(n229), .IN5(n3508), 
        .IN6(n197), .Q(n1276) );
  NAND4X0 U389 ( .IN1(n1283), .IN2(n1284), .IN3(n1285), .IN4(n1286), .QN(n1274) );
  OA221X1 U390 ( .IN1(n3505), .IN2(n101), .IN3(n3502), .IN4(n69), .IN5(n1287), 
        .Q(n1286) );
  OA22X1 U391 ( .IN1(n3499), .IN2(n133), .IN3(n3496), .IN4(n37), .Q(n1287) );
  OA221X1 U392 ( .IN1(n3493), .IN2(n901), .IN3(n3490), .IN4(n933), .IN5(n1288), 
        .Q(n1285) );
  OA22X1 U393 ( .IN1(n3487), .IN2(n5), .IN3(n3484), .IN4(n965), .Q(n1288) );
  OA221X1 U394 ( .IN1(n3481), .IN2(n773), .IN3(n3478), .IN4(n805), .IN5(n1289), 
        .Q(n1284) );
  OA22X1 U395 ( .IN1(n3475), .IN2(n869), .IN3(n3472), .IN4(n837), .Q(n1289) );
  OA221X1 U396 ( .IN1(n3469), .IN2(n709), .IN3(n3466), .IN4(n741), .IN5(n1290), 
        .Q(n1283) );
  OA22X1 U397 ( .IN1(n3463), .IN2(n677), .IN3(n3460), .IN4(n645), .Q(n1290) );
  OR2X1 U398 ( .IN1(n1291), .IN2(n1292), .Q(rd_dataB[26]) );
  NAND4X0 U399 ( .IN1(n1293), .IN2(n1294), .IN3(n1295), .IN4(n1296), .QN(n1292) );
  OA221X1 U400 ( .IN1(n3550), .IN2(n518), .IN3(n3547), .IN4(n550), .IN5(n1297), 
        .Q(n1296) );
  OA22X1 U401 ( .IN1(n3544), .IN2(n614), .IN3(n3541), .IN4(n582), .Q(n1297) );
  OA221X1 U402 ( .IN1(n3538), .IN2(n390), .IN3(n3535), .IN4(n422), .IN5(n1298), 
        .Q(n1295) );
  OA22X1 U403 ( .IN1(n3532), .IN2(n486), .IN3(n3529), .IN4(n454), .Q(n1298) );
  OA221X1 U404 ( .IN1(n3526), .IN2(n262), .IN3(n3523), .IN4(n294), .IN5(n1299), 
        .Q(n1294) );
  OA22X1 U405 ( .IN1(n3520), .IN2(n358), .IN3(n3517), .IN4(n326), .Q(n1299) );
  OA222X1 U406 ( .IN1(n3514), .IN2(n166), .IN3(n3511), .IN4(n230), .IN5(n3508), 
        .IN6(n198), .Q(n1293) );
  NAND4X0 U407 ( .IN1(n1300), .IN2(n1301), .IN3(n1302), .IN4(n1303), .QN(n1291) );
  OA221X1 U408 ( .IN1(n3505), .IN2(n102), .IN3(n3502), .IN4(n70), .IN5(n1304), 
        .Q(n1303) );
  OA22X1 U409 ( .IN1(n3499), .IN2(n134), .IN3(n3496), .IN4(n38), .Q(n1304) );
  OA221X1 U410 ( .IN1(n3493), .IN2(n902), .IN3(n3490), .IN4(n934), .IN5(n1305), 
        .Q(n1302) );
  OA22X1 U411 ( .IN1(n3487), .IN2(n6), .IN3(n3484), .IN4(n966), .Q(n1305) );
  OA221X1 U412 ( .IN1(n3481), .IN2(n774), .IN3(n3478), .IN4(n806), .IN5(n1306), 
        .Q(n1301) );
  OA22X1 U413 ( .IN1(n3475), .IN2(n870), .IN3(n3472), .IN4(n838), .Q(n1306) );
  OA221X1 U414 ( .IN1(n3469), .IN2(n710), .IN3(n3466), .IN4(n742), .IN5(n1307), 
        .Q(n1300) );
  OA22X1 U415 ( .IN1(n3463), .IN2(n678), .IN3(n3460), .IN4(n646), .Q(n1307) );
  OR2X1 U416 ( .IN1(n1308), .IN2(n1309), .Q(rd_dataB[25]) );
  NAND4X0 U417 ( .IN1(n1310), .IN2(n1311), .IN3(n1312), .IN4(n1313), .QN(n1309) );
  OA221X1 U418 ( .IN1(n3550), .IN2(n519), .IN3(n3547), .IN4(n551), .IN5(n1314), 
        .Q(n1313) );
  OA22X1 U419 ( .IN1(n3544), .IN2(n615), .IN3(n3541), .IN4(n583), .Q(n1314) );
  OA221X1 U420 ( .IN1(n3538), .IN2(n391), .IN3(n3535), .IN4(n423), .IN5(n1315), 
        .Q(n1312) );
  OA22X1 U421 ( .IN1(n3532), .IN2(n487), .IN3(n3529), .IN4(n455), .Q(n1315) );
  OA221X1 U422 ( .IN1(n3526), .IN2(n263), .IN3(n3523), .IN4(n295), .IN5(n1316), 
        .Q(n1311) );
  OA22X1 U423 ( .IN1(n3520), .IN2(n359), .IN3(n3517), .IN4(n327), .Q(n1316) );
  OA222X1 U424 ( .IN1(n3514), .IN2(n167), .IN3(n3511), .IN4(n231), .IN5(n3508), 
        .IN6(n199), .Q(n1310) );
  NAND4X0 U425 ( .IN1(n1317), .IN2(n1318), .IN3(n1319), .IN4(n1320), .QN(n1308) );
  OA221X1 U426 ( .IN1(n3505), .IN2(n103), .IN3(n3502), .IN4(n71), .IN5(n1321), 
        .Q(n1320) );
  OA22X1 U427 ( .IN1(n3499), .IN2(n135), .IN3(n3496), .IN4(n39), .Q(n1321) );
  OA221X1 U428 ( .IN1(n3493), .IN2(n903), .IN3(n3490), .IN4(n935), .IN5(n1322), 
        .Q(n1319) );
  OA22X1 U429 ( .IN1(n3487), .IN2(n7), .IN3(n3484), .IN4(n967), .Q(n1322) );
  OA221X1 U430 ( .IN1(n3481), .IN2(n775), .IN3(n3478), .IN4(n807), .IN5(n1323), 
        .Q(n1318) );
  OA22X1 U431 ( .IN1(n3475), .IN2(n871), .IN3(n3472), .IN4(n839), .Q(n1323) );
  OA221X1 U432 ( .IN1(n3469), .IN2(n711), .IN3(n3466), .IN4(n743), .IN5(n1324), 
        .Q(n1317) );
  OA22X1 U433 ( .IN1(n3463), .IN2(n679), .IN3(n3460), .IN4(n647), .Q(n1324) );
  OR2X1 U434 ( .IN1(n1325), .IN2(n1326), .Q(rd_dataB[24]) );
  NAND4X0 U435 ( .IN1(n1327), .IN2(n1328), .IN3(n1329), .IN4(n1330), .QN(n1326) );
  OA221X1 U436 ( .IN1(n3550), .IN2(n520), .IN3(n3547), .IN4(n552), .IN5(n1331), 
        .Q(n1330) );
  OA22X1 U437 ( .IN1(n3544), .IN2(n616), .IN3(n3541), .IN4(n584), .Q(n1331) );
  OA221X1 U438 ( .IN1(n3538), .IN2(n392), .IN3(n3535), .IN4(n424), .IN5(n1332), 
        .Q(n1329) );
  OA22X1 U439 ( .IN1(n3532), .IN2(n488), .IN3(n3529), .IN4(n456), .Q(n1332) );
  OA221X1 U440 ( .IN1(n3526), .IN2(n264), .IN3(n3523), .IN4(n296), .IN5(n1333), 
        .Q(n1328) );
  OA22X1 U441 ( .IN1(n3520), .IN2(n360), .IN3(n3517), .IN4(n328), .Q(n1333) );
  OA222X1 U442 ( .IN1(n3514), .IN2(n168), .IN3(n3511), .IN4(n232), .IN5(n3508), 
        .IN6(n200), .Q(n1327) );
  NAND4X0 U443 ( .IN1(n1334), .IN2(n1335), .IN3(n1336), .IN4(n1337), .QN(n1325) );
  OA221X1 U444 ( .IN1(n3505), .IN2(n104), .IN3(n3502), .IN4(n72), .IN5(n1338), 
        .Q(n1337) );
  OA22X1 U445 ( .IN1(n3499), .IN2(n136), .IN3(n3496), .IN4(n40), .Q(n1338) );
  OA221X1 U446 ( .IN1(n3493), .IN2(n904), .IN3(n3490), .IN4(n936), .IN5(n1339), 
        .Q(n1336) );
  OA22X1 U447 ( .IN1(n3487), .IN2(n8), .IN3(n3484), .IN4(n968), .Q(n1339) );
  OA221X1 U448 ( .IN1(n3481), .IN2(n776), .IN3(n3478), .IN4(n808), .IN5(n1340), 
        .Q(n1335) );
  OA22X1 U449 ( .IN1(n3475), .IN2(n872), .IN3(n3472), .IN4(n840), .Q(n1340) );
  OA221X1 U450 ( .IN1(n3469), .IN2(n712), .IN3(n3466), .IN4(n744), .IN5(n1341), 
        .Q(n1334) );
  OA22X1 U451 ( .IN1(n3463), .IN2(n680), .IN3(n3460), .IN4(n648), .Q(n1341) );
  OR2X1 U452 ( .IN1(n1342), .IN2(n1343), .Q(rd_dataB[23]) );
  NAND4X0 U453 ( .IN1(n1344), .IN2(n1345), .IN3(n1346), .IN4(n1347), .QN(n1343) );
  OA221X1 U454 ( .IN1(n3550), .IN2(n521), .IN3(n3547), .IN4(n553), .IN5(n1348), 
        .Q(n1347) );
  OA22X1 U455 ( .IN1(n3544), .IN2(n617), .IN3(n3541), .IN4(n585), .Q(n1348) );
  OA221X1 U456 ( .IN1(n3538), .IN2(n393), .IN3(n3535), .IN4(n425), .IN5(n1349), 
        .Q(n1346) );
  OA22X1 U457 ( .IN1(n3532), .IN2(n489), .IN3(n3529), .IN4(n457), .Q(n1349) );
  OA221X1 U458 ( .IN1(n3526), .IN2(n265), .IN3(n3523), .IN4(n297), .IN5(n1350), 
        .Q(n1345) );
  OA22X1 U459 ( .IN1(n3520), .IN2(n361), .IN3(n3517), .IN4(n329), .Q(n1350) );
  OA222X1 U460 ( .IN1(n3514), .IN2(n169), .IN3(n3511), .IN4(n233), .IN5(n3508), 
        .IN6(n201), .Q(n1344) );
  NAND4X0 U461 ( .IN1(n1351), .IN2(n1352), .IN3(n1353), .IN4(n1354), .QN(n1342) );
  OA221X1 U462 ( .IN1(n3505), .IN2(n105), .IN3(n3502), .IN4(n73), .IN5(n1355), 
        .Q(n1354) );
  OA22X1 U463 ( .IN1(n3499), .IN2(n137), .IN3(n3496), .IN4(n41), .Q(n1355) );
  OA221X1 U464 ( .IN1(n3493), .IN2(n905), .IN3(n3490), .IN4(n937), .IN5(n1356), 
        .Q(n1353) );
  OA22X1 U465 ( .IN1(n3487), .IN2(n9), .IN3(n3484), .IN4(n969), .Q(n1356) );
  OA221X1 U466 ( .IN1(n3481), .IN2(n777), .IN3(n3478), .IN4(n809), .IN5(n1357), 
        .Q(n1352) );
  OA22X1 U467 ( .IN1(n3475), .IN2(n873), .IN3(n3472), .IN4(n841), .Q(n1357) );
  OA221X1 U468 ( .IN1(n3469), .IN2(n713), .IN3(n3466), .IN4(n745), .IN5(n1358), 
        .Q(n1351) );
  OA22X1 U469 ( .IN1(n3463), .IN2(n681), .IN3(n3460), .IN4(n649), .Q(n1358) );
  OR2X1 U470 ( .IN1(n1359), .IN2(n1360), .Q(rd_dataB[22]) );
  NAND4X0 U471 ( .IN1(n1361), .IN2(n1362), .IN3(n1363), .IN4(n1364), .QN(n1360) );
  OA221X1 U472 ( .IN1(n3550), .IN2(n522), .IN3(n3547), .IN4(n554), .IN5(n1365), 
        .Q(n1364) );
  OA22X1 U473 ( .IN1(n3544), .IN2(n618), .IN3(n3541), .IN4(n586), .Q(n1365) );
  OA221X1 U474 ( .IN1(n3538), .IN2(n394), .IN3(n3535), .IN4(n426), .IN5(n1366), 
        .Q(n1363) );
  OA22X1 U475 ( .IN1(n3532), .IN2(n490), .IN3(n3529), .IN4(n458), .Q(n1366) );
  OA221X1 U476 ( .IN1(n3526), .IN2(n266), .IN3(n3523), .IN4(n298), .IN5(n1367), 
        .Q(n1362) );
  OA22X1 U477 ( .IN1(n3520), .IN2(n362), .IN3(n3517), .IN4(n330), .Q(n1367) );
  OA222X1 U478 ( .IN1(n3514), .IN2(n170), .IN3(n3511), .IN4(n234), .IN5(n3508), 
        .IN6(n202), .Q(n1361) );
  NAND4X0 U479 ( .IN1(n1368), .IN2(n1369), .IN3(n1370), .IN4(n1371), .QN(n1359) );
  OA221X1 U480 ( .IN1(n3505), .IN2(n106), .IN3(n3502), .IN4(n74), .IN5(n1372), 
        .Q(n1371) );
  OA22X1 U481 ( .IN1(n3499), .IN2(n138), .IN3(n3496), .IN4(n42), .Q(n1372) );
  OA221X1 U482 ( .IN1(n3493), .IN2(n906), .IN3(n3490), .IN4(n938), .IN5(n1373), 
        .Q(n1370) );
  OA22X1 U483 ( .IN1(n3487), .IN2(n10), .IN3(n3484), .IN4(n970), .Q(n1373) );
  OA221X1 U484 ( .IN1(n3481), .IN2(n778), .IN3(n3478), .IN4(n810), .IN5(n1374), 
        .Q(n1369) );
  OA22X1 U485 ( .IN1(n3475), .IN2(n874), .IN3(n3472), .IN4(n842), .Q(n1374) );
  OA221X1 U486 ( .IN1(n3469), .IN2(n714), .IN3(n3466), .IN4(n746), .IN5(n1375), 
        .Q(n1368) );
  OA22X1 U487 ( .IN1(n3463), .IN2(n682), .IN3(n3460), .IN4(n650), .Q(n1375) );
  OR2X1 U488 ( .IN1(n1376), .IN2(n1377), .Q(rd_dataB[21]) );
  NAND4X0 U489 ( .IN1(n1378), .IN2(n1379), .IN3(n1380), .IN4(n1381), .QN(n1377) );
  OA221X1 U490 ( .IN1(n3550), .IN2(n523), .IN3(n3547), .IN4(n555), .IN5(n1382), 
        .Q(n1381) );
  OA22X1 U491 ( .IN1(n3544), .IN2(n619), .IN3(n3541), .IN4(n587), .Q(n1382) );
  OA221X1 U492 ( .IN1(n3538), .IN2(n395), .IN3(n3535), .IN4(n427), .IN5(n1383), 
        .Q(n1380) );
  OA22X1 U493 ( .IN1(n3532), .IN2(n491), .IN3(n3529), .IN4(n459), .Q(n1383) );
  OA221X1 U494 ( .IN1(n3526), .IN2(n267), .IN3(n3523), .IN4(n299), .IN5(n1384), 
        .Q(n1379) );
  OA22X1 U495 ( .IN1(n3520), .IN2(n363), .IN3(n3517), .IN4(n331), .Q(n1384) );
  OA222X1 U496 ( .IN1(n3514), .IN2(n171), .IN3(n3511), .IN4(n235), .IN5(n3508), 
        .IN6(n203), .Q(n1378) );
  NAND4X0 U497 ( .IN1(n1385), .IN2(n1386), .IN3(n1387), .IN4(n1388), .QN(n1376) );
  OA221X1 U498 ( .IN1(n3505), .IN2(n107), .IN3(n3502), .IN4(n75), .IN5(n1389), 
        .Q(n1388) );
  OA22X1 U499 ( .IN1(n3499), .IN2(n139), .IN3(n3496), .IN4(n43), .Q(n1389) );
  OA221X1 U500 ( .IN1(n3493), .IN2(n907), .IN3(n3490), .IN4(n939), .IN5(n1390), 
        .Q(n1387) );
  OA22X1 U501 ( .IN1(n3487), .IN2(n11), .IN3(n3484), .IN4(n971), .Q(n1390) );
  OA221X1 U502 ( .IN1(n3481), .IN2(n779), .IN3(n3478), .IN4(n811), .IN5(n1391), 
        .Q(n1386) );
  OA22X1 U503 ( .IN1(n3475), .IN2(n875), .IN3(n3472), .IN4(n843), .Q(n1391) );
  OA221X1 U504 ( .IN1(n3469), .IN2(n715), .IN3(n3466), .IN4(n747), .IN5(n1392), 
        .Q(n1385) );
  OA22X1 U505 ( .IN1(n3463), .IN2(n683), .IN3(n3460), .IN4(n651), .Q(n1392) );
  OR2X1 U506 ( .IN1(n1393), .IN2(n1394), .Q(rd_dataB[20]) );
  NAND4X0 U507 ( .IN1(n1395), .IN2(n1396), .IN3(n1397), .IN4(n1398), .QN(n1394) );
  OA221X1 U508 ( .IN1(n3550), .IN2(n524), .IN3(n3547), .IN4(n556), .IN5(n1399), 
        .Q(n1398) );
  OA22X1 U509 ( .IN1(n3544), .IN2(n620), .IN3(n3541), .IN4(n588), .Q(n1399) );
  OA221X1 U510 ( .IN1(n3538), .IN2(n396), .IN3(n3535), .IN4(n428), .IN5(n1400), 
        .Q(n1397) );
  OA22X1 U511 ( .IN1(n3532), .IN2(n492), .IN3(n3529), .IN4(n460), .Q(n1400) );
  OA221X1 U512 ( .IN1(n3526), .IN2(n268), .IN3(n3523), .IN4(n300), .IN5(n1401), 
        .Q(n1396) );
  OA22X1 U513 ( .IN1(n3520), .IN2(n364), .IN3(n3517), .IN4(n332), .Q(n1401) );
  OA222X1 U514 ( .IN1(n3514), .IN2(n172), .IN3(n3511), .IN4(n236), .IN5(n3508), 
        .IN6(n204), .Q(n1395) );
  NAND4X0 U515 ( .IN1(n1402), .IN2(n1403), .IN3(n1404), .IN4(n1405), .QN(n1393) );
  OA221X1 U516 ( .IN1(n3505), .IN2(n108), .IN3(n3502), .IN4(n76), .IN5(n1406), 
        .Q(n1405) );
  OA22X1 U517 ( .IN1(n3499), .IN2(n140), .IN3(n3496), .IN4(n44), .Q(n1406) );
  OA221X1 U518 ( .IN1(n3493), .IN2(n908), .IN3(n3490), .IN4(n940), .IN5(n1407), 
        .Q(n1404) );
  OA22X1 U519 ( .IN1(n3487), .IN2(n12), .IN3(n3484), .IN4(n972), .Q(n1407) );
  OA221X1 U520 ( .IN1(n3481), .IN2(n780), .IN3(n3478), .IN4(n812), .IN5(n1408), 
        .Q(n1403) );
  OA22X1 U521 ( .IN1(n3475), .IN2(n876), .IN3(n3472), .IN4(n844), .Q(n1408) );
  OA221X1 U522 ( .IN1(n3469), .IN2(n716), .IN3(n3466), .IN4(n748), .IN5(n1409), 
        .Q(n1402) );
  OA22X1 U523 ( .IN1(n3463), .IN2(n684), .IN3(n3460), .IN4(n652), .Q(n1409) );
  OR2X1 U524 ( .IN1(n1410), .IN2(n1411), .Q(rd_dataB[1]) );
  NAND4X0 U525 ( .IN1(n1412), .IN2(n1413), .IN3(n1414), .IN4(n1415), .QN(n1411) );
  OA221X1 U526 ( .IN1(n3550), .IN2(n543), .IN3(n3547), .IN4(n575), .IN5(n1416), 
        .Q(n1415) );
  OA22X1 U527 ( .IN1(n3544), .IN2(n639), .IN3(n3541), .IN4(n607), .Q(n1416) );
  OA221X1 U528 ( .IN1(n3538), .IN2(n415), .IN3(n3535), .IN4(n447), .IN5(n1417), 
        .Q(n1414) );
  OA22X1 U529 ( .IN1(n3532), .IN2(n511), .IN3(n3529), .IN4(n479), .Q(n1417) );
  OA221X1 U530 ( .IN1(n3526), .IN2(n287), .IN3(n3523), .IN4(n319), .IN5(n1418), 
        .Q(n1413) );
  OA22X1 U531 ( .IN1(n3520), .IN2(n383), .IN3(n3517), .IN4(n351), .Q(n1418) );
  OA222X1 U532 ( .IN1(n3514), .IN2(n191), .IN3(n3511), .IN4(n255), .IN5(n3508), 
        .IN6(n223), .Q(n1412) );
  NAND4X0 U533 ( .IN1(n1419), .IN2(n1420), .IN3(n1421), .IN4(n1422), .QN(n1410) );
  OA221X1 U534 ( .IN1(n3505), .IN2(n127), .IN3(n3502), .IN4(n95), .IN5(n1423), 
        .Q(n1422) );
  OA22X1 U535 ( .IN1(n3499), .IN2(n159), .IN3(n3496), .IN4(n63), .Q(n1423) );
  OA221X1 U536 ( .IN1(n3493), .IN2(n927), .IN3(n3490), .IN4(n959), .IN5(n1424), 
        .Q(n1421) );
  OA22X1 U537 ( .IN1(n3487), .IN2(n31), .IN3(n3484), .IN4(n991), .Q(n1424) );
  OA221X1 U538 ( .IN1(n3481), .IN2(n799), .IN3(n3478), .IN4(n831), .IN5(n1425), 
        .Q(n1420) );
  OA22X1 U539 ( .IN1(n3475), .IN2(n895), .IN3(n3472), .IN4(n863), .Q(n1425) );
  OA221X1 U540 ( .IN1(n3469), .IN2(n735), .IN3(n3466), .IN4(n767), .IN5(n1426), 
        .Q(n1419) );
  OA22X1 U541 ( .IN1(n3463), .IN2(n703), .IN3(n3460), .IN4(n671), .Q(n1426) );
  OR2X1 U542 ( .IN1(n1427), .IN2(n1428), .Q(rd_dataB[19]) );
  NAND4X0 U543 ( .IN1(n1429), .IN2(n1430), .IN3(n1431), .IN4(n1432), .QN(n1428) );
  OA221X1 U544 ( .IN1(n3550), .IN2(n525), .IN3(n3547), .IN4(n557), .IN5(n1433), 
        .Q(n1432) );
  OA22X1 U545 ( .IN1(n3544), .IN2(n621), .IN3(n3541), .IN4(n589), .Q(n1433) );
  OA221X1 U546 ( .IN1(n3538), .IN2(n397), .IN3(n3535), .IN4(n429), .IN5(n1434), 
        .Q(n1431) );
  OA22X1 U547 ( .IN1(n3532), .IN2(n493), .IN3(n3529), .IN4(n461), .Q(n1434) );
  OA221X1 U548 ( .IN1(n3526), .IN2(n269), .IN3(n3523), .IN4(n301), .IN5(n1435), 
        .Q(n1430) );
  OA22X1 U549 ( .IN1(n3520), .IN2(n365), .IN3(n3517), .IN4(n333), .Q(n1435) );
  OA222X1 U550 ( .IN1(n3514), .IN2(n173), .IN3(n3511), .IN4(n237), .IN5(n3508), 
        .IN6(n205), .Q(n1429) );
  NAND4X0 U551 ( .IN1(n1436), .IN2(n1437), .IN3(n1438), .IN4(n1439), .QN(n1427) );
  OA221X1 U552 ( .IN1(n3505), .IN2(n109), .IN3(n3502), .IN4(n77), .IN5(n1440), 
        .Q(n1439) );
  OA22X1 U553 ( .IN1(n3499), .IN2(n141), .IN3(n3496), .IN4(n45), .Q(n1440) );
  OA221X1 U554 ( .IN1(n3493), .IN2(n909), .IN3(n3490), .IN4(n941), .IN5(n1441), 
        .Q(n1438) );
  OA22X1 U555 ( .IN1(n3487), .IN2(n13), .IN3(n3484), .IN4(n973), .Q(n1441) );
  OA221X1 U556 ( .IN1(n3481), .IN2(n781), .IN3(n3478), .IN4(n813), .IN5(n1442), 
        .Q(n1437) );
  OA22X1 U557 ( .IN1(n3475), .IN2(n877), .IN3(n3472), .IN4(n845), .Q(n1442) );
  OA221X1 U558 ( .IN1(n3469), .IN2(n717), .IN3(n3466), .IN4(n749), .IN5(n1443), 
        .Q(n1436) );
  OA22X1 U559 ( .IN1(n3463), .IN2(n685), .IN3(n3460), .IN4(n653), .Q(n1443) );
  OR2X1 U560 ( .IN1(n1444), .IN2(n1445), .Q(rd_dataB[18]) );
  NAND4X0 U561 ( .IN1(n1446), .IN2(n1447), .IN3(n1448), .IN4(n1449), .QN(n1445) );
  OA221X1 U562 ( .IN1(n3550), .IN2(n526), .IN3(n3547), .IN4(n558), .IN5(n1450), 
        .Q(n1449) );
  OA22X1 U563 ( .IN1(n3544), .IN2(n622), .IN3(n3541), .IN4(n590), .Q(n1450) );
  OA221X1 U564 ( .IN1(n3538), .IN2(n398), .IN3(n3535), .IN4(n430), .IN5(n1451), 
        .Q(n1448) );
  OA22X1 U565 ( .IN1(n3532), .IN2(n494), .IN3(n3529), .IN4(n462), .Q(n1451) );
  OA221X1 U566 ( .IN1(n3526), .IN2(n270), .IN3(n3523), .IN4(n302), .IN5(n1452), 
        .Q(n1447) );
  OA22X1 U567 ( .IN1(n3520), .IN2(n366), .IN3(n3517), .IN4(n334), .Q(n1452) );
  OA222X1 U568 ( .IN1(n3514), .IN2(n174), .IN3(n3511), .IN4(n238), .IN5(n3508), 
        .IN6(n206), .Q(n1446) );
  NAND4X0 U569 ( .IN1(n1453), .IN2(n1454), .IN3(n1455), .IN4(n1456), .QN(n1444) );
  OA221X1 U570 ( .IN1(n3505), .IN2(n110), .IN3(n3502), .IN4(n78), .IN5(n1457), 
        .Q(n1456) );
  OA22X1 U571 ( .IN1(n3499), .IN2(n142), .IN3(n3496), .IN4(n46), .Q(n1457) );
  OA221X1 U572 ( .IN1(n3493), .IN2(n910), .IN3(n3490), .IN4(n942), .IN5(n1458), 
        .Q(n1455) );
  OA22X1 U573 ( .IN1(n3487), .IN2(n14), .IN3(n3484), .IN4(n974), .Q(n1458) );
  OA221X1 U574 ( .IN1(n3481), .IN2(n782), .IN3(n3478), .IN4(n814), .IN5(n1459), 
        .Q(n1454) );
  OA22X1 U575 ( .IN1(n3475), .IN2(n878), .IN3(n3472), .IN4(n846), .Q(n1459) );
  OA221X1 U576 ( .IN1(n3469), .IN2(n718), .IN3(n3466), .IN4(n750), .IN5(n1460), 
        .Q(n1453) );
  OA22X1 U577 ( .IN1(n3463), .IN2(n686), .IN3(n3460), .IN4(n654), .Q(n1460) );
  OR2X1 U578 ( .IN1(n1461), .IN2(n1462), .Q(rd_dataB[17]) );
  NAND4X0 U579 ( .IN1(n1463), .IN2(n1464), .IN3(n1465), .IN4(n1466), .QN(n1462) );
  OA221X1 U580 ( .IN1(n3550), .IN2(n527), .IN3(n3547), .IN4(n559), .IN5(n1467), 
        .Q(n1466) );
  OA22X1 U581 ( .IN1(n3544), .IN2(n623), .IN3(n3541), .IN4(n591), .Q(n1467) );
  OA221X1 U582 ( .IN1(n3538), .IN2(n399), .IN3(n3535), .IN4(n431), .IN5(n1468), 
        .Q(n1465) );
  OA22X1 U583 ( .IN1(n3532), .IN2(n495), .IN3(n3529), .IN4(n463), .Q(n1468) );
  OA221X1 U584 ( .IN1(n3526), .IN2(n271), .IN3(n3523), .IN4(n303), .IN5(n1469), 
        .Q(n1464) );
  OA22X1 U585 ( .IN1(n3520), .IN2(n367), .IN3(n3517), .IN4(n335), .Q(n1469) );
  OA222X1 U586 ( .IN1(n3514), .IN2(n175), .IN3(n3511), .IN4(n239), .IN5(n3508), 
        .IN6(n207), .Q(n1463) );
  NAND4X0 U587 ( .IN1(n1470), .IN2(n1471), .IN3(n1472), .IN4(n1473), .QN(n1461) );
  OA221X1 U588 ( .IN1(n3505), .IN2(n111), .IN3(n3502), .IN4(n79), .IN5(n1474), 
        .Q(n1473) );
  OA22X1 U589 ( .IN1(n3499), .IN2(n143), .IN3(n3496), .IN4(n47), .Q(n1474) );
  OA221X1 U590 ( .IN1(n3493), .IN2(n911), .IN3(n3490), .IN4(n943), .IN5(n1475), 
        .Q(n1472) );
  OA22X1 U591 ( .IN1(n3487), .IN2(n15), .IN3(n3484), .IN4(n975), .Q(n1475) );
  OA221X1 U592 ( .IN1(n3481), .IN2(n783), .IN3(n3478), .IN4(n815), .IN5(n1476), 
        .Q(n1471) );
  OA22X1 U593 ( .IN1(n3475), .IN2(n879), .IN3(n3472), .IN4(n847), .Q(n1476) );
  OA221X1 U594 ( .IN1(n3469), .IN2(n719), .IN3(n3466), .IN4(n751), .IN5(n1477), 
        .Q(n1470) );
  OA22X1 U595 ( .IN1(n3463), .IN2(n687), .IN3(n3460), .IN4(n655), .Q(n1477) );
  OR2X1 U596 ( .IN1(n1478), .IN2(n1479), .Q(rd_dataB[16]) );
  NAND4X0 U597 ( .IN1(n1480), .IN2(n1481), .IN3(n1482), .IN4(n1483), .QN(n1479) );
  OA221X1 U598 ( .IN1(n3551), .IN2(n528), .IN3(n3548), .IN4(n560), .IN5(n1484), 
        .Q(n1483) );
  OA22X1 U599 ( .IN1(n3545), .IN2(n624), .IN3(n3542), .IN4(n592), .Q(n1484) );
  OA221X1 U600 ( .IN1(n3539), .IN2(n400), .IN3(n3536), .IN4(n432), .IN5(n1485), 
        .Q(n1482) );
  OA22X1 U601 ( .IN1(n3533), .IN2(n496), .IN3(n3530), .IN4(n464), .Q(n1485) );
  OA221X1 U602 ( .IN1(n3527), .IN2(n272), .IN3(n3524), .IN4(n304), .IN5(n1486), 
        .Q(n1481) );
  OA22X1 U603 ( .IN1(n3521), .IN2(n368), .IN3(n3518), .IN4(n336), .Q(n1486) );
  OA222X1 U604 ( .IN1(n3515), .IN2(n176), .IN3(n3512), .IN4(n240), .IN5(n3509), 
        .IN6(n208), .Q(n1480) );
  NAND4X0 U605 ( .IN1(n1487), .IN2(n1488), .IN3(n1489), .IN4(n1490), .QN(n1478) );
  OA221X1 U606 ( .IN1(n3506), .IN2(n112), .IN3(n3503), .IN4(n80), .IN5(n1491), 
        .Q(n1490) );
  OA22X1 U607 ( .IN1(n3500), .IN2(n144), .IN3(n3497), .IN4(n48), .Q(n1491) );
  OA221X1 U608 ( .IN1(n3494), .IN2(n912), .IN3(n3491), .IN4(n944), .IN5(n1492), 
        .Q(n1489) );
  OA22X1 U609 ( .IN1(n3488), .IN2(n16), .IN3(n3485), .IN4(n976), .Q(n1492) );
  OA221X1 U610 ( .IN1(n3482), .IN2(n784), .IN3(n3479), .IN4(n816), .IN5(n1493), 
        .Q(n1488) );
  OA22X1 U611 ( .IN1(n3476), .IN2(n880), .IN3(n3473), .IN4(n848), .Q(n1493) );
  OA221X1 U612 ( .IN1(n3470), .IN2(n720), .IN3(n3467), .IN4(n752), .IN5(n1494), 
        .Q(n1487) );
  OA22X1 U613 ( .IN1(n3464), .IN2(n688), .IN3(n3461), .IN4(n656), .Q(n1494) );
  OR2X1 U614 ( .IN1(n1495), .IN2(n1496), .Q(rd_dataB[15]) );
  NAND4X0 U615 ( .IN1(n1497), .IN2(n1498), .IN3(n1499), .IN4(n1500), .QN(n1496) );
  OA221X1 U616 ( .IN1(n3551), .IN2(n529), .IN3(n3548), .IN4(n561), .IN5(n1501), 
        .Q(n1500) );
  OA22X1 U617 ( .IN1(n3545), .IN2(n625), .IN3(n3542), .IN4(n593), .Q(n1501) );
  OA221X1 U618 ( .IN1(n3539), .IN2(n401), .IN3(n3536), .IN4(n433), .IN5(n1502), 
        .Q(n1499) );
  OA22X1 U619 ( .IN1(n3533), .IN2(n497), .IN3(n3530), .IN4(n465), .Q(n1502) );
  OA221X1 U620 ( .IN1(n3527), .IN2(n273), .IN3(n3524), .IN4(n305), .IN5(n1503), 
        .Q(n1498) );
  OA22X1 U621 ( .IN1(n3521), .IN2(n369), .IN3(n3518), .IN4(n337), .Q(n1503) );
  OA222X1 U622 ( .IN1(n3515), .IN2(n177), .IN3(n3512), .IN4(n241), .IN5(n3509), 
        .IN6(n209), .Q(n1497) );
  NAND4X0 U623 ( .IN1(n1504), .IN2(n1505), .IN3(n1506), .IN4(n1507), .QN(n1495) );
  OA221X1 U624 ( .IN1(n3506), .IN2(n113), .IN3(n3503), .IN4(n81), .IN5(n1508), 
        .Q(n1507) );
  OA22X1 U625 ( .IN1(n3500), .IN2(n145), .IN3(n3497), .IN4(n49), .Q(n1508) );
  OA221X1 U626 ( .IN1(n3494), .IN2(n913), .IN3(n3491), .IN4(n945), .IN5(n1509), 
        .Q(n1506) );
  OA22X1 U627 ( .IN1(n3488), .IN2(n17), .IN3(n3485), .IN4(n977), .Q(n1509) );
  OA221X1 U628 ( .IN1(n3482), .IN2(n785), .IN3(n3479), .IN4(n817), .IN5(n1510), 
        .Q(n1505) );
  OA22X1 U629 ( .IN1(n3476), .IN2(n881), .IN3(n3473), .IN4(n849), .Q(n1510) );
  OA221X1 U630 ( .IN1(n3470), .IN2(n721), .IN3(n3467), .IN4(n753), .IN5(n1511), 
        .Q(n1504) );
  OA22X1 U631 ( .IN1(n3464), .IN2(n689), .IN3(n3461), .IN4(n657), .Q(n1511) );
  OR2X1 U632 ( .IN1(n1512), .IN2(n1513), .Q(rd_dataB[14]) );
  NAND4X0 U633 ( .IN1(n1514), .IN2(n1515), .IN3(n1516), .IN4(n1517), .QN(n1513) );
  OA221X1 U634 ( .IN1(n3551), .IN2(n530), .IN3(n3548), .IN4(n562), .IN5(n1518), 
        .Q(n1517) );
  OA22X1 U635 ( .IN1(n3545), .IN2(n626), .IN3(n3542), .IN4(n594), .Q(n1518) );
  OA221X1 U636 ( .IN1(n3539), .IN2(n402), .IN3(n3536), .IN4(n434), .IN5(n1519), 
        .Q(n1516) );
  OA22X1 U637 ( .IN1(n3533), .IN2(n498), .IN3(n3530), .IN4(n466), .Q(n1519) );
  OA221X1 U638 ( .IN1(n3527), .IN2(n274), .IN3(n3524), .IN4(n306), .IN5(n1520), 
        .Q(n1515) );
  OA22X1 U639 ( .IN1(n3521), .IN2(n370), .IN3(n3518), .IN4(n338), .Q(n1520) );
  OA222X1 U640 ( .IN1(n3515), .IN2(n178), .IN3(n3512), .IN4(n242), .IN5(n3509), 
        .IN6(n210), .Q(n1514) );
  NAND4X0 U641 ( .IN1(n1521), .IN2(n1522), .IN3(n1523), .IN4(n1524), .QN(n1512) );
  OA221X1 U642 ( .IN1(n3506), .IN2(n114), .IN3(n3503), .IN4(n82), .IN5(n1525), 
        .Q(n1524) );
  OA22X1 U643 ( .IN1(n3500), .IN2(n146), .IN3(n3497), .IN4(n50), .Q(n1525) );
  OA221X1 U644 ( .IN1(n3494), .IN2(n914), .IN3(n3491), .IN4(n946), .IN5(n1526), 
        .Q(n1523) );
  OA22X1 U645 ( .IN1(n3488), .IN2(n18), .IN3(n3485), .IN4(n978), .Q(n1526) );
  OA221X1 U646 ( .IN1(n3482), .IN2(n786), .IN3(n3479), .IN4(n818), .IN5(n1527), 
        .Q(n1522) );
  OA22X1 U647 ( .IN1(n3476), .IN2(n882), .IN3(n3473), .IN4(n850), .Q(n1527) );
  OA221X1 U648 ( .IN1(n3470), .IN2(n722), .IN3(n3467), .IN4(n754), .IN5(n1528), 
        .Q(n1521) );
  OA22X1 U649 ( .IN1(n3464), .IN2(n690), .IN3(n3461), .IN4(n658), .Q(n1528) );
  OR2X1 U650 ( .IN1(n1529), .IN2(n1530), .Q(rd_dataB[13]) );
  NAND4X0 U651 ( .IN1(n1531), .IN2(n1532), .IN3(n1533), .IN4(n1534), .QN(n1530) );
  OA221X1 U652 ( .IN1(n3551), .IN2(n531), .IN3(n3548), .IN4(n563), .IN5(n1535), 
        .Q(n1534) );
  OA22X1 U653 ( .IN1(n3545), .IN2(n627), .IN3(n3542), .IN4(n595), .Q(n1535) );
  OA221X1 U654 ( .IN1(n3539), .IN2(n403), .IN3(n3536), .IN4(n435), .IN5(n1536), 
        .Q(n1533) );
  OA22X1 U655 ( .IN1(n3533), .IN2(n499), .IN3(n3530), .IN4(n467), .Q(n1536) );
  OA221X1 U656 ( .IN1(n3527), .IN2(n275), .IN3(n3524), .IN4(n307), .IN5(n1537), 
        .Q(n1532) );
  OA22X1 U657 ( .IN1(n3521), .IN2(n371), .IN3(n3518), .IN4(n339), .Q(n1537) );
  OA222X1 U658 ( .IN1(n3515), .IN2(n179), .IN3(n3512), .IN4(n243), .IN5(n3509), 
        .IN6(n211), .Q(n1531) );
  NAND4X0 U659 ( .IN1(n1538), .IN2(n1539), .IN3(n1540), .IN4(n1541), .QN(n1529) );
  OA221X1 U660 ( .IN1(n3506), .IN2(n115), .IN3(n3503), .IN4(n83), .IN5(n1542), 
        .Q(n1541) );
  OA22X1 U661 ( .IN1(n3500), .IN2(n147), .IN3(n3497), .IN4(n51), .Q(n1542) );
  OA221X1 U662 ( .IN1(n3494), .IN2(n915), .IN3(n3491), .IN4(n947), .IN5(n1543), 
        .Q(n1540) );
  OA22X1 U663 ( .IN1(n3488), .IN2(n19), .IN3(n3485), .IN4(n979), .Q(n1543) );
  OA221X1 U664 ( .IN1(n3482), .IN2(n787), .IN3(n3479), .IN4(n819), .IN5(n1544), 
        .Q(n1539) );
  OA22X1 U665 ( .IN1(n3476), .IN2(n883), .IN3(n3473), .IN4(n851), .Q(n1544) );
  OA221X1 U666 ( .IN1(n3470), .IN2(n723), .IN3(n3467), .IN4(n755), .IN5(n1545), 
        .Q(n1538) );
  OA22X1 U667 ( .IN1(n3464), .IN2(n691), .IN3(n3461), .IN4(n659), .Q(n1545) );
  OR2X1 U668 ( .IN1(n1546), .IN2(n1547), .Q(rd_dataB[12]) );
  NAND4X0 U669 ( .IN1(n1548), .IN2(n1549), .IN3(n1550), .IN4(n1551), .QN(n1547) );
  OA221X1 U670 ( .IN1(n3551), .IN2(n532), .IN3(n3548), .IN4(n564), .IN5(n1552), 
        .Q(n1551) );
  OA22X1 U671 ( .IN1(n3545), .IN2(n628), .IN3(n3542), .IN4(n596), .Q(n1552) );
  OA221X1 U672 ( .IN1(n3539), .IN2(n404), .IN3(n3536), .IN4(n436), .IN5(n1553), 
        .Q(n1550) );
  OA22X1 U673 ( .IN1(n3533), .IN2(n500), .IN3(n3530), .IN4(n468), .Q(n1553) );
  OA221X1 U674 ( .IN1(n3527), .IN2(n276), .IN3(n3524), .IN4(n308), .IN5(n1554), 
        .Q(n1549) );
  OA22X1 U675 ( .IN1(n3521), .IN2(n372), .IN3(n3518), .IN4(n340), .Q(n1554) );
  OA222X1 U676 ( .IN1(n3515), .IN2(n180), .IN3(n3512), .IN4(n244), .IN5(n3509), 
        .IN6(n212), .Q(n1548) );
  NAND4X0 U677 ( .IN1(n1555), .IN2(n1556), .IN3(n1557), .IN4(n1558), .QN(n1546) );
  OA221X1 U678 ( .IN1(n3506), .IN2(n116), .IN3(n3503), .IN4(n84), .IN5(n1559), 
        .Q(n1558) );
  OA22X1 U679 ( .IN1(n3500), .IN2(n148), .IN3(n3497), .IN4(n52), .Q(n1559) );
  OA221X1 U680 ( .IN1(n3494), .IN2(n916), .IN3(n3491), .IN4(n948), .IN5(n1560), 
        .Q(n1557) );
  OA22X1 U681 ( .IN1(n3488), .IN2(n20), .IN3(n3485), .IN4(n980), .Q(n1560) );
  OA221X1 U682 ( .IN1(n3482), .IN2(n788), .IN3(n3479), .IN4(n820), .IN5(n1561), 
        .Q(n1556) );
  OA22X1 U683 ( .IN1(n3476), .IN2(n884), .IN3(n3473), .IN4(n852), .Q(n1561) );
  OA221X1 U684 ( .IN1(n3470), .IN2(n724), .IN3(n3467), .IN4(n756), .IN5(n1562), 
        .Q(n1555) );
  OA22X1 U685 ( .IN1(n3464), .IN2(n692), .IN3(n3461), .IN4(n660), .Q(n1562) );
  OR2X1 U686 ( .IN1(n1563), .IN2(n1564), .Q(rd_dataB[11]) );
  NAND4X0 U687 ( .IN1(n1565), .IN2(n1566), .IN3(n1567), .IN4(n1568), .QN(n1564) );
  OA221X1 U688 ( .IN1(n3551), .IN2(n533), .IN3(n3548), .IN4(n565), .IN5(n1569), 
        .Q(n1568) );
  OA22X1 U689 ( .IN1(n3545), .IN2(n629), .IN3(n3542), .IN4(n597), .Q(n1569) );
  OA221X1 U690 ( .IN1(n3539), .IN2(n405), .IN3(n3536), .IN4(n437), .IN5(n1570), 
        .Q(n1567) );
  OA22X1 U691 ( .IN1(n3533), .IN2(n501), .IN3(n3530), .IN4(n469), .Q(n1570) );
  OA221X1 U692 ( .IN1(n3527), .IN2(n277), .IN3(n3524), .IN4(n309), .IN5(n1571), 
        .Q(n1566) );
  OA22X1 U693 ( .IN1(n3521), .IN2(n373), .IN3(n3518), .IN4(n341), .Q(n1571) );
  OA222X1 U694 ( .IN1(n3515), .IN2(n181), .IN3(n3512), .IN4(n245), .IN5(n3509), 
        .IN6(n213), .Q(n1565) );
  NAND4X0 U695 ( .IN1(n1572), .IN2(n1573), .IN3(n1574), .IN4(n1575), .QN(n1563) );
  OA221X1 U696 ( .IN1(n3506), .IN2(n117), .IN3(n3503), .IN4(n85), .IN5(n1576), 
        .Q(n1575) );
  OA22X1 U697 ( .IN1(n3500), .IN2(n149), .IN3(n3497), .IN4(n53), .Q(n1576) );
  OA221X1 U698 ( .IN1(n3494), .IN2(n917), .IN3(n3491), .IN4(n949), .IN5(n1577), 
        .Q(n1574) );
  OA22X1 U699 ( .IN1(n3488), .IN2(n21), .IN3(n3485), .IN4(n981), .Q(n1577) );
  OA221X1 U700 ( .IN1(n3482), .IN2(n789), .IN3(n3479), .IN4(n821), .IN5(n1578), 
        .Q(n1573) );
  OA22X1 U701 ( .IN1(n3476), .IN2(n885), .IN3(n3473), .IN4(n853), .Q(n1578) );
  OA221X1 U702 ( .IN1(n3470), .IN2(n725), .IN3(n3467), .IN4(n757), .IN5(n1579), 
        .Q(n1572) );
  OA22X1 U703 ( .IN1(n3464), .IN2(n693), .IN3(n3461), .IN4(n661), .Q(n1579) );
  OR2X1 U704 ( .IN1(n1580), .IN2(n1581), .Q(rd_dataB[10]) );
  NAND4X0 U705 ( .IN1(n1582), .IN2(n1583), .IN3(n1584), .IN4(n1585), .QN(n1581) );
  OA221X1 U706 ( .IN1(n3551), .IN2(n534), .IN3(n3548), .IN4(n566), .IN5(n1586), 
        .Q(n1585) );
  OA22X1 U707 ( .IN1(n3545), .IN2(n630), .IN3(n3542), .IN4(n598), .Q(n1586) );
  OA221X1 U708 ( .IN1(n3539), .IN2(n406), .IN3(n3536), .IN4(n438), .IN5(n1587), 
        .Q(n1584) );
  OA22X1 U709 ( .IN1(n3533), .IN2(n502), .IN3(n3530), .IN4(n470), .Q(n1587) );
  OA221X1 U710 ( .IN1(n3527), .IN2(n278), .IN3(n3524), .IN4(n310), .IN5(n1588), 
        .Q(n1583) );
  OA22X1 U711 ( .IN1(n3521), .IN2(n374), .IN3(n3518), .IN4(n342), .Q(n1588) );
  OA222X1 U712 ( .IN1(n3515), .IN2(n182), .IN3(n3512), .IN4(n246), .IN5(n3509), 
        .IN6(n214), .Q(n1582) );
  NAND4X0 U713 ( .IN1(n1589), .IN2(n1590), .IN3(n1591), .IN4(n1592), .QN(n1580) );
  OA221X1 U714 ( .IN1(n3506), .IN2(n118), .IN3(n3503), .IN4(n86), .IN5(n1593), 
        .Q(n1592) );
  OA22X1 U715 ( .IN1(n3500), .IN2(n150), .IN3(n3497), .IN4(n54), .Q(n1593) );
  OA221X1 U716 ( .IN1(n3494), .IN2(n918), .IN3(n3491), .IN4(n950), .IN5(n1594), 
        .Q(n1591) );
  OA22X1 U717 ( .IN1(n3488), .IN2(n22), .IN3(n3485), .IN4(n982), .Q(n1594) );
  OA221X1 U718 ( .IN1(n3482), .IN2(n790), .IN3(n3479), .IN4(n822), .IN5(n1595), 
        .Q(n1590) );
  OA22X1 U719 ( .IN1(n3476), .IN2(n886), .IN3(n3473), .IN4(n854), .Q(n1595) );
  OA221X1 U720 ( .IN1(n3470), .IN2(n726), .IN3(n3467), .IN4(n758), .IN5(n1596), 
        .Q(n1589) );
  OA22X1 U721 ( .IN1(n3464), .IN2(n694), .IN3(n3461), .IN4(n662), .Q(n1596) );
  OR2X1 U722 ( .IN1(n1597), .IN2(n1598), .Q(rd_dataB[0]) );
  NAND4X0 U723 ( .IN1(n1599), .IN2(n1600), .IN3(n1601), .IN4(n1602), .QN(n1598) );
  OA221X1 U724 ( .IN1(n3551), .IN2(n544), .IN3(n3548), .IN4(n576), .IN5(n1603), 
        .Q(n1602) );
  OA22X1 U725 ( .IN1(n3545), .IN2(n640), .IN3(n3542), .IN4(n608), .Q(n1603) );
  OA221X1 U726 ( .IN1(n3539), .IN2(n416), .IN3(n3536), .IN4(n448), .IN5(n1608), 
        .Q(n1601) );
  OA22X1 U727 ( .IN1(n3533), .IN2(n512), .IN3(n3530), .IN4(n480), .Q(n1608) );
  OA221X1 U728 ( .IN1(n3527), .IN2(n288), .IN3(n3524), .IN4(n320), .IN5(n1611), 
        .Q(n1600) );
  OA22X1 U729 ( .IN1(n3521), .IN2(n384), .IN3(n3518), .IN4(n352), .Q(n1611) );
  OA222X1 U730 ( .IN1(n3515), .IN2(n192), .IN3(n3512), .IN4(n256), .IN5(n3509), 
        .IN6(n224), .Q(n1599) );
  NAND4X0 U731 ( .IN1(n1616), .IN2(n1617), .IN3(n1618), .IN4(n1619), .QN(n1597) );
  OA221X1 U732 ( .IN1(n3506), .IN2(n128), .IN3(n3503), .IN4(n96), .IN5(n1620), 
        .Q(n1619) );
  OA22X1 U733 ( .IN1(n3500), .IN2(n160), .IN3(n3497), .IN4(n64), .Q(n1620) );
  AND3X1 U734 ( .IN1(rd_addrB[2]), .IN2(rd_addrB[1]), .IN3(rd_addrB[3]), .Q(
        n1605) );
  AND2X1 U735 ( .IN1(n1623), .IN2(rd_addrB[3]), .Q(n1607) );
  OA221X1 U736 ( .IN1(n3494), .IN2(n928), .IN3(n3491), .IN4(n960), .IN5(n1624), 
        .Q(n1618) );
  OA22X1 U737 ( .IN1(n3488), .IN2(n32), .IN3(n3485), .IN4(n992), .Q(n1624) );
  AND2X1 U738 ( .IN1(n1625), .IN2(rd_addrB[1]), .Q(n1609) );
  AND2X1 U739 ( .IN1(n1625), .IN2(n3751), .Q(n1610) );
  OA221X1 U740 ( .IN1(n3482), .IN2(n800), .IN3(n3479), .IN4(n832), .IN5(n1626), 
        .Q(n1617) );
  OA22X1 U741 ( .IN1(n3476), .IN2(n896), .IN3(n3473), .IN4(n864), .Q(n1626) );
  AND2X1 U742 ( .IN1(n1627), .IN2(rd_addrB[2]), .Q(n1612) );
  AND2X1 U743 ( .IN1(n1623), .IN2(n3749), .Q(n1613) );
  OA221X1 U744 ( .IN1(n3470), .IN2(n736), .IN3(n3467), .IN4(n768), .IN5(n1628), 
        .Q(n1616) );
  OA22X1 U745 ( .IN1(n3464), .IN2(n704), .IN3(n3461), .IN4(n672), .Q(n1628) );
  AND3X1 U746 ( .IN1(n3750), .IN2(n3749), .IN3(n3751), .Q(n1615) );
  AND2X1 U747 ( .IN1(n1627), .IN2(n3750), .Q(n1614) );
  OR2X1 U748 ( .IN1(n1629), .IN2(n1630), .Q(rd_dataA[9]) );
  NAND4X0 U749 ( .IN1(n1631), .IN2(n1632), .IN3(n1633), .IN4(n1634), .QN(n1630) );
  OA221X1 U750 ( .IN1(n535), .IN2(n3456), .IN3(n567), .IN4(n3453), .IN5(n1637), 
        .Q(n1634) );
  OA22X1 U751 ( .IN1(n631), .IN2(n3450), .IN3(n599), .IN4(n3447), .Q(n1637) );
  OA221X1 U752 ( .IN1(n407), .IN2(n3444), .IN3(n439), .IN4(n3441), .IN5(n1642), 
        .Q(n1633) );
  OA22X1 U753 ( .IN1(n503), .IN2(n3438), .IN3(n471), .IN4(n3435), .Q(n1642) );
  OA221X1 U754 ( .IN1(n279), .IN2(n3432), .IN3(n311), .IN4(n3429), .IN5(n1647), 
        .Q(n1632) );
  OA22X1 U755 ( .IN1(n375), .IN2(n3426), .IN3(n343), .IN4(n3423), .Q(n1647) );
  OA222X1 U756 ( .IN1(n183), .IN2(n3420), .IN3(n247), .IN4(n3417), .IN5(n215), 
        .IN6(n3414), .Q(n1631) );
  NAND4X0 U757 ( .IN1(n1653), .IN2(n1654), .IN3(n1655), .IN4(n1656), .QN(n1629) );
  OA221X1 U758 ( .IN1(n119), .IN2(n3411), .IN3(n87), .IN4(n3408), .IN5(n1659), 
        .Q(n1656) );
  OA22X1 U759 ( .IN1(n151), .IN2(n3405), .IN3(n55), .IN4(n3402), .Q(n1659) );
  OA221X1 U760 ( .IN1(n919), .IN2(n3399), .IN3(n951), .IN4(n3396), .IN5(n1664), 
        .Q(n1655) );
  OA22X1 U761 ( .IN1(n23), .IN2(n3393), .IN3(n983), .IN4(n3390), .Q(n1664) );
  OA221X1 U762 ( .IN1(n791), .IN2(n3387), .IN3(n823), .IN4(n3384), .IN5(n1669), 
        .Q(n1654) );
  OA22X1 U763 ( .IN1(n887), .IN2(n3381), .IN3(n855), .IN4(n3378), .Q(n1669) );
  OA221X1 U764 ( .IN1(n727), .IN2(n3375), .IN3(n759), .IN4(n3372), .IN5(n1674), 
        .Q(n1653) );
  OA22X1 U765 ( .IN1(n695), .IN2(n3369), .IN3(n663), .IN4(n3366), .Q(n1674) );
  OR2X1 U766 ( .IN1(n1677), .IN2(n1678), .Q(rd_dataA[8]) );
  NAND4X0 U767 ( .IN1(n1679), .IN2(n1680), .IN3(n1681), .IN4(n1682), .QN(n1678) );
  OA221X1 U768 ( .IN1(n536), .IN2(n3456), .IN3(n568), .IN4(n3453), .IN5(n1683), 
        .Q(n1682) );
  OA22X1 U769 ( .IN1(n632), .IN2(n3450), .IN3(n600), .IN4(n3447), .Q(n1683) );
  OA221X1 U770 ( .IN1(n408), .IN2(n3444), .IN3(n440), .IN4(n3441), .IN5(n1684), 
        .Q(n1681) );
  OA22X1 U771 ( .IN1(n504), .IN2(n3438), .IN3(n472), .IN4(n3435), .Q(n1684) );
  OA221X1 U772 ( .IN1(n280), .IN2(n3432), .IN3(n312), .IN4(n3429), .IN5(n1685), 
        .Q(n1680) );
  OA22X1 U773 ( .IN1(n376), .IN2(n3426), .IN3(n344), .IN4(n3423), .Q(n1685) );
  OA222X1 U774 ( .IN1(n184), .IN2(n3420), .IN3(n248), .IN4(n3417), .IN5(n216), 
        .IN6(n3414), .Q(n1679) );
  NAND4X0 U775 ( .IN1(n1686), .IN2(n1687), .IN3(n1688), .IN4(n1689), .QN(n1677) );
  OA221X1 U776 ( .IN1(n120), .IN2(n3411), .IN3(n88), .IN4(n3408), .IN5(n1690), 
        .Q(n1689) );
  OA22X1 U777 ( .IN1(n152), .IN2(n3405), .IN3(n56), .IN4(n3402), .Q(n1690) );
  OA221X1 U778 ( .IN1(n920), .IN2(n3399), .IN3(n952), .IN4(n3396), .IN5(n1691), 
        .Q(n1688) );
  OA22X1 U779 ( .IN1(n24), .IN2(n3393), .IN3(n984), .IN4(n3390), .Q(n1691) );
  OA221X1 U780 ( .IN1(n792), .IN2(n3387), .IN3(n824), .IN4(n3384), .IN5(n1692), 
        .Q(n1687) );
  OA22X1 U781 ( .IN1(n888), .IN2(n3381), .IN3(n856), .IN4(n3378), .Q(n1692) );
  OA221X1 U782 ( .IN1(n728), .IN2(n3375), .IN3(n760), .IN4(n3372), .IN5(n1693), 
        .Q(n1686) );
  OA22X1 U783 ( .IN1(n696), .IN2(n3369), .IN3(n664), .IN4(n3366), .Q(n1693) );
  OR2X1 U784 ( .IN1(n1694), .IN2(n1695), .Q(rd_dataA[7]) );
  NAND4X0 U785 ( .IN1(n1696), .IN2(n1697), .IN3(n1698), .IN4(n1699), .QN(n1695) );
  OA221X1 U786 ( .IN1(n537), .IN2(n3456), .IN3(n569), .IN4(n3453), .IN5(n1700), 
        .Q(n1699) );
  OA22X1 U787 ( .IN1(n633), .IN2(n3450), .IN3(n601), .IN4(n3447), .Q(n1700) );
  OA221X1 U788 ( .IN1(n409), .IN2(n3444), .IN3(n441), .IN4(n3441), .IN5(n1701), 
        .Q(n1698) );
  OA22X1 U789 ( .IN1(n505), .IN2(n3438), .IN3(n473), .IN4(n3435), .Q(n1701) );
  OA221X1 U790 ( .IN1(n281), .IN2(n3432), .IN3(n313), .IN4(n3429), .IN5(n1702), 
        .Q(n1697) );
  OA22X1 U791 ( .IN1(n377), .IN2(n3426), .IN3(n345), .IN4(n3423), .Q(n1702) );
  OA222X1 U792 ( .IN1(n185), .IN2(n3420), .IN3(n249), .IN4(n3417), .IN5(n217), 
        .IN6(n3414), .Q(n1696) );
  NAND4X0 U793 ( .IN1(n1703), .IN2(n1704), .IN3(n1705), .IN4(n1706), .QN(n1694) );
  OA221X1 U794 ( .IN1(n121), .IN2(n3411), .IN3(n89), .IN4(n3408), .IN5(n1707), 
        .Q(n1706) );
  OA22X1 U795 ( .IN1(n153), .IN2(n3405), .IN3(n57), .IN4(n3402), .Q(n1707) );
  OA221X1 U796 ( .IN1(n921), .IN2(n3399), .IN3(n953), .IN4(n3396), .IN5(n1708), 
        .Q(n1705) );
  OA22X1 U797 ( .IN1(n25), .IN2(n3393), .IN3(n985), .IN4(n3390), .Q(n1708) );
  OA221X1 U798 ( .IN1(n793), .IN2(n3387), .IN3(n825), .IN4(n3384), .IN5(n1709), 
        .Q(n1704) );
  OA22X1 U799 ( .IN1(n889), .IN2(n3381), .IN3(n857), .IN4(n3378), .Q(n1709) );
  OA221X1 U800 ( .IN1(n729), .IN2(n3375), .IN3(n761), .IN4(n3372), .IN5(n1710), 
        .Q(n1703) );
  OA22X1 U801 ( .IN1(n697), .IN2(n3369), .IN3(n665), .IN4(n3366), .Q(n1710) );
  OR2X1 U802 ( .IN1(n1711), .IN2(n1712), .Q(rd_dataA[6]) );
  NAND4X0 U803 ( .IN1(n1713), .IN2(n1714), .IN3(n1715), .IN4(n1716), .QN(n1712) );
  OA221X1 U804 ( .IN1(n538), .IN2(n3456), .IN3(n570), .IN4(n3453), .IN5(n1717), 
        .Q(n1716) );
  OA22X1 U805 ( .IN1(n634), .IN2(n3450), .IN3(n602), .IN4(n3447), .Q(n1717) );
  OA221X1 U806 ( .IN1(n410), .IN2(n3444), .IN3(n442), .IN4(n3441), .IN5(n1718), 
        .Q(n1715) );
  OA22X1 U807 ( .IN1(n506), .IN2(n3438), .IN3(n474), .IN4(n3435), .Q(n1718) );
  OA221X1 U808 ( .IN1(n282), .IN2(n3432), .IN3(n314), .IN4(n3429), .IN5(n1719), 
        .Q(n1714) );
  OA22X1 U809 ( .IN1(n378), .IN2(n3426), .IN3(n346), .IN4(n3423), .Q(n1719) );
  OA222X1 U810 ( .IN1(n186), .IN2(n3420), .IN3(n250), .IN4(n3417), .IN5(n218), 
        .IN6(n3414), .Q(n1713) );
  NAND4X0 U811 ( .IN1(n1720), .IN2(n1721), .IN3(n1722), .IN4(n1723), .QN(n1711) );
  OA221X1 U812 ( .IN1(n122), .IN2(n3411), .IN3(n90), .IN4(n3408), .IN5(n1724), 
        .Q(n1723) );
  OA22X1 U813 ( .IN1(n154), .IN2(n3405), .IN3(n58), .IN4(n3402), .Q(n1724) );
  OA221X1 U814 ( .IN1(n922), .IN2(n3399), .IN3(n954), .IN4(n3396), .IN5(n1725), 
        .Q(n1722) );
  OA22X1 U815 ( .IN1(n26), .IN2(n3393), .IN3(n986), .IN4(n3390), .Q(n1725) );
  OA221X1 U816 ( .IN1(n794), .IN2(n3387), .IN3(n826), .IN4(n3384), .IN5(n1726), 
        .Q(n1721) );
  OA22X1 U817 ( .IN1(n890), .IN2(n3381), .IN3(n858), .IN4(n3378), .Q(n1726) );
  OA221X1 U818 ( .IN1(n730), .IN2(n3375), .IN3(n762), .IN4(n3372), .IN5(n1727), 
        .Q(n1720) );
  OA22X1 U819 ( .IN1(n698), .IN2(n3369), .IN3(n666), .IN4(n3366), .Q(n1727) );
  OR2X1 U820 ( .IN1(n1728), .IN2(n1729), .Q(rd_dataA[5]) );
  NAND4X0 U821 ( .IN1(n1730), .IN2(n1731), .IN3(n1732), .IN4(n1733), .QN(n1729) );
  OA221X1 U822 ( .IN1(n539), .IN2(n3456), .IN3(n571), .IN4(n3453), .IN5(n1734), 
        .Q(n1733) );
  OA22X1 U823 ( .IN1(n635), .IN2(n3450), .IN3(n603), .IN4(n3447), .Q(n1734) );
  OA221X1 U824 ( .IN1(n411), .IN2(n3444), .IN3(n443), .IN4(n3441), .IN5(n1735), 
        .Q(n1732) );
  OA22X1 U825 ( .IN1(n507), .IN2(n3438), .IN3(n475), .IN4(n3435), .Q(n1735) );
  OA221X1 U826 ( .IN1(n283), .IN2(n3432), .IN3(n315), .IN4(n3429), .IN5(n1736), 
        .Q(n1731) );
  OA22X1 U827 ( .IN1(n379), .IN2(n3426), .IN3(n347), .IN4(n3423), .Q(n1736) );
  OA222X1 U828 ( .IN1(n187), .IN2(n3420), .IN3(n251), .IN4(n3417), .IN5(n219), 
        .IN6(n3414), .Q(n1730) );
  NAND4X0 U829 ( .IN1(n1737), .IN2(n1738), .IN3(n1739), .IN4(n1740), .QN(n1728) );
  OA221X1 U830 ( .IN1(n123), .IN2(n3411), .IN3(n91), .IN4(n3408), .IN5(n1741), 
        .Q(n1740) );
  OA22X1 U831 ( .IN1(n155), .IN2(n3405), .IN3(n59), .IN4(n3402), .Q(n1741) );
  OA221X1 U832 ( .IN1(n923), .IN2(n3399), .IN3(n955), .IN4(n3396), .IN5(n1742), 
        .Q(n1739) );
  OA22X1 U833 ( .IN1(n27), .IN2(n3393), .IN3(n987), .IN4(n3390), .Q(n1742) );
  OA221X1 U834 ( .IN1(n795), .IN2(n3387), .IN3(n827), .IN4(n3384), .IN5(n1743), 
        .Q(n1738) );
  OA22X1 U835 ( .IN1(n891), .IN2(n3381), .IN3(n859), .IN4(n3378), .Q(n1743) );
  OA221X1 U836 ( .IN1(n731), .IN2(n3375), .IN3(n763), .IN4(n3372), .IN5(n1744), 
        .Q(n1737) );
  OA22X1 U837 ( .IN1(n699), .IN2(n3369), .IN3(n667), .IN4(n3366), .Q(n1744) );
  OR2X1 U838 ( .IN1(n1745), .IN2(n1746), .Q(rd_dataA[4]) );
  NAND4X0 U839 ( .IN1(n1747), .IN2(n1748), .IN3(n1749), .IN4(n1750), .QN(n1746) );
  OA221X1 U840 ( .IN1(n540), .IN2(n3456), .IN3(n572), .IN4(n3453), .IN5(n1751), 
        .Q(n1750) );
  OA22X1 U841 ( .IN1(n636), .IN2(n3450), .IN3(n604), .IN4(n3447), .Q(n1751) );
  OA221X1 U842 ( .IN1(n412), .IN2(n3444), .IN3(n444), .IN4(n3441), .IN5(n1752), 
        .Q(n1749) );
  OA22X1 U843 ( .IN1(n508), .IN2(n3438), .IN3(n476), .IN4(n3435), .Q(n1752) );
  OA221X1 U844 ( .IN1(n284), .IN2(n3432), .IN3(n316), .IN4(n3429), .IN5(n1753), 
        .Q(n1748) );
  OA22X1 U845 ( .IN1(n380), .IN2(n3426), .IN3(n348), .IN4(n3423), .Q(n1753) );
  OA222X1 U846 ( .IN1(n188), .IN2(n3420), .IN3(n252), .IN4(n3417), .IN5(n220), 
        .IN6(n3414), .Q(n1747) );
  NAND4X0 U847 ( .IN1(n1754), .IN2(n1755), .IN3(n1756), .IN4(n1757), .QN(n1745) );
  OA221X1 U848 ( .IN1(n124), .IN2(n3411), .IN3(n92), .IN4(n3408), .IN5(n1758), 
        .Q(n1757) );
  OA22X1 U849 ( .IN1(n156), .IN2(n3405), .IN3(n60), .IN4(n3402), .Q(n1758) );
  OA221X1 U850 ( .IN1(n924), .IN2(n3399), .IN3(n956), .IN4(n3396), .IN5(n1759), 
        .Q(n1756) );
  OA22X1 U851 ( .IN1(n28), .IN2(n3393), .IN3(n988), .IN4(n3390), .Q(n1759) );
  OA221X1 U852 ( .IN1(n796), .IN2(n3387), .IN3(n828), .IN4(n3384), .IN5(n1760), 
        .Q(n1755) );
  OA22X1 U853 ( .IN1(n892), .IN2(n3381), .IN3(n860), .IN4(n3378), .Q(n1760) );
  OA221X1 U854 ( .IN1(n732), .IN2(n3375), .IN3(n764), .IN4(n3372), .IN5(n1761), 
        .Q(n1754) );
  OA22X1 U855 ( .IN1(n700), .IN2(n3369), .IN3(n668), .IN4(n3366), .Q(n1761) );
  OR2X1 U856 ( .IN1(n1762), .IN2(n1763), .Q(rd_dataA[3]) );
  NAND4X0 U857 ( .IN1(n1764), .IN2(n1765), .IN3(n1766), .IN4(n1767), .QN(n1763) );
  OA221X1 U858 ( .IN1(n541), .IN2(n3456), .IN3(n573), .IN4(n3453), .IN5(n1768), 
        .Q(n1767) );
  OA22X1 U859 ( .IN1(n637), .IN2(n3450), .IN3(n605), .IN4(n3447), .Q(n1768) );
  OA221X1 U860 ( .IN1(n413), .IN2(n3444), .IN3(n445), .IN4(n3441), .IN5(n1769), 
        .Q(n1766) );
  OA22X1 U861 ( .IN1(n509), .IN2(n3438), .IN3(n477), .IN4(n3435), .Q(n1769) );
  OA221X1 U862 ( .IN1(n285), .IN2(n3432), .IN3(n317), .IN4(n3429), .IN5(n1770), 
        .Q(n1765) );
  OA22X1 U863 ( .IN1(n381), .IN2(n3426), .IN3(n349), .IN4(n3423), .Q(n1770) );
  OA222X1 U864 ( .IN1(n189), .IN2(n3420), .IN3(n253), .IN4(n3417), .IN5(n221), 
        .IN6(n3414), .Q(n1764) );
  NAND4X0 U865 ( .IN1(n1771), .IN2(n1772), .IN3(n1773), .IN4(n1774), .QN(n1762) );
  OA221X1 U866 ( .IN1(n125), .IN2(n3411), .IN3(n93), .IN4(n3408), .IN5(n1775), 
        .Q(n1774) );
  OA22X1 U867 ( .IN1(n157), .IN2(n3405), .IN3(n61), .IN4(n3402), .Q(n1775) );
  OA221X1 U868 ( .IN1(n925), .IN2(n3399), .IN3(n957), .IN4(n3396), .IN5(n1776), 
        .Q(n1773) );
  OA22X1 U869 ( .IN1(n29), .IN2(n3393), .IN3(n989), .IN4(n3390), .Q(n1776) );
  OA221X1 U870 ( .IN1(n797), .IN2(n3387), .IN3(n829), .IN4(n3384), .IN5(n1777), 
        .Q(n1772) );
  OA22X1 U871 ( .IN1(n893), .IN2(n3381), .IN3(n861), .IN4(n3378), .Q(n1777) );
  OA221X1 U872 ( .IN1(n733), .IN2(n3375), .IN3(n765), .IN4(n3372), .IN5(n1778), 
        .Q(n1771) );
  OA22X1 U873 ( .IN1(n701), .IN2(n3369), .IN3(n669), .IN4(n3366), .Q(n1778) );
  OR2X1 U874 ( .IN1(n1779), .IN2(n1780), .Q(rd_dataA[31]) );
  NAND4X0 U875 ( .IN1(n1781), .IN2(n1782), .IN3(n1783), .IN4(n1784), .QN(n1780) );
  OA221X1 U876 ( .IN1(n513), .IN2(n3456), .IN3(n545), .IN4(n3453), .IN5(n1785), 
        .Q(n1784) );
  OA22X1 U877 ( .IN1(n609), .IN2(n3450), .IN3(n577), .IN4(n3447), .Q(n1785) );
  OA221X1 U878 ( .IN1(n385), .IN2(n3444), .IN3(n417), .IN4(n3441), .IN5(n1786), 
        .Q(n1783) );
  OA22X1 U879 ( .IN1(n481), .IN2(n3438), .IN3(n449), .IN4(n3435), .Q(n1786) );
  OA221X1 U880 ( .IN1(n257), .IN2(n3432), .IN3(n289), .IN4(n3429), .IN5(n1787), 
        .Q(n1782) );
  OA22X1 U881 ( .IN1(n353), .IN2(n3426), .IN3(n321), .IN4(n3423), .Q(n1787) );
  OA222X1 U882 ( .IN1(n161), .IN2(n3420), .IN3(n225), .IN4(n3417), .IN5(n193), 
        .IN6(n3414), .Q(n1781) );
  NAND4X0 U883 ( .IN1(n1788), .IN2(n1789), .IN3(n1790), .IN4(n1791), .QN(n1779) );
  OA221X1 U884 ( .IN1(n97), .IN2(n3411), .IN3(n65), .IN4(n3408), .IN5(n1792), 
        .Q(n1791) );
  OA22X1 U885 ( .IN1(n129), .IN2(n3405), .IN3(n33), .IN4(n3402), .Q(n1792) );
  OA221X1 U886 ( .IN1(n897), .IN2(n3399), .IN3(n929), .IN4(n3396), .IN5(n1793), 
        .Q(n1790) );
  OA22X1 U887 ( .IN1(n1), .IN2(n3393), .IN3(n961), .IN4(n3390), .Q(n1793) );
  OA221X1 U888 ( .IN1(n769), .IN2(n3387), .IN3(n801), .IN4(n3384), .IN5(n1794), 
        .Q(n1789) );
  OA22X1 U889 ( .IN1(n865), .IN2(n3381), .IN3(n833), .IN4(n3378), .Q(n1794) );
  OA221X1 U890 ( .IN1(n705), .IN2(n3375), .IN3(n737), .IN4(n3372), .IN5(n1795), 
        .Q(n1788) );
  OA22X1 U891 ( .IN1(n673), .IN2(n3369), .IN3(n641), .IN4(n3366), .Q(n1795) );
  OR2X1 U892 ( .IN1(n1796), .IN2(n1797), .Q(rd_dataA[30]) );
  NAND4X0 U893 ( .IN1(n1798), .IN2(n1799), .IN3(n1800), .IN4(n1801), .QN(n1797) );
  OA221X1 U894 ( .IN1(n514), .IN2(n3456), .IN3(n546), .IN4(n3453), .IN5(n1802), 
        .Q(n1801) );
  OA22X1 U895 ( .IN1(n610), .IN2(n3450), .IN3(n578), .IN4(n3447), .Q(n1802) );
  OA221X1 U896 ( .IN1(n386), .IN2(n3444), .IN3(n418), .IN4(n3441), .IN5(n1803), 
        .Q(n1800) );
  OA22X1 U897 ( .IN1(n482), .IN2(n3438), .IN3(n450), .IN4(n3435), .Q(n1803) );
  OA221X1 U898 ( .IN1(n258), .IN2(n3432), .IN3(n290), .IN4(n3429), .IN5(n1804), 
        .Q(n1799) );
  OA22X1 U899 ( .IN1(n354), .IN2(n3426), .IN3(n322), .IN4(n3423), .Q(n1804) );
  OA222X1 U900 ( .IN1(n162), .IN2(n3420), .IN3(n226), .IN4(n3417), .IN5(n194), 
        .IN6(n3414), .Q(n1798) );
  NAND4X0 U901 ( .IN1(n1805), .IN2(n1806), .IN3(n1807), .IN4(n1808), .QN(n1796) );
  OA221X1 U902 ( .IN1(n98), .IN2(n3411), .IN3(n66), .IN4(n3408), .IN5(n1809), 
        .Q(n1808) );
  OA22X1 U903 ( .IN1(n130), .IN2(n3405), .IN3(n34), .IN4(n3402), .Q(n1809) );
  OA221X1 U904 ( .IN1(n898), .IN2(n3399), .IN3(n930), .IN4(n3396), .IN5(n1810), 
        .Q(n1807) );
  OA22X1 U905 ( .IN1(n2), .IN2(n3393), .IN3(n962), .IN4(n3390), .Q(n1810) );
  OA221X1 U906 ( .IN1(n770), .IN2(n3387), .IN3(n802), .IN4(n3384), .IN5(n1811), 
        .Q(n1806) );
  OA22X1 U907 ( .IN1(n866), .IN2(n3381), .IN3(n834), .IN4(n3378), .Q(n1811) );
  OA221X1 U908 ( .IN1(n706), .IN2(n3375), .IN3(n738), .IN4(n3372), .IN5(n1812), 
        .Q(n1805) );
  OA22X1 U909 ( .IN1(n674), .IN2(n3369), .IN3(n642), .IN4(n3366), .Q(n1812) );
  OR2X1 U910 ( .IN1(n1813), .IN2(n1814), .Q(rd_dataA[2]) );
  NAND4X0 U911 ( .IN1(n1815), .IN2(n1816), .IN3(n1817), .IN4(n1818), .QN(n1814) );
  OA221X1 U912 ( .IN1(n542), .IN2(n3456), .IN3(n574), .IN4(n3453), .IN5(n1819), 
        .Q(n1818) );
  OA22X1 U913 ( .IN1(n638), .IN2(n3450), .IN3(n606), .IN4(n3447), .Q(n1819) );
  OA221X1 U914 ( .IN1(n414), .IN2(n3444), .IN3(n446), .IN4(n3441), .IN5(n1820), 
        .Q(n1817) );
  OA22X1 U915 ( .IN1(n510), .IN2(n3438), .IN3(n478), .IN4(n3435), .Q(n1820) );
  OA221X1 U916 ( .IN1(n286), .IN2(n3432), .IN3(n318), .IN4(n3429), .IN5(n1821), 
        .Q(n1816) );
  OA22X1 U917 ( .IN1(n382), .IN2(n3426), .IN3(n350), .IN4(n3423), .Q(n1821) );
  OA222X1 U918 ( .IN1(n190), .IN2(n3420), .IN3(n254), .IN4(n3417), .IN5(n222), 
        .IN6(n3414), .Q(n1815) );
  NAND4X0 U919 ( .IN1(n1822), .IN2(n1823), .IN3(n1824), .IN4(n1825), .QN(n1813) );
  OA221X1 U920 ( .IN1(n126), .IN2(n3411), .IN3(n94), .IN4(n3408), .IN5(n1826), 
        .Q(n1825) );
  OA22X1 U921 ( .IN1(n158), .IN2(n3405), .IN3(n62), .IN4(n3402), .Q(n1826) );
  OA221X1 U922 ( .IN1(n926), .IN2(n3399), .IN3(n958), .IN4(n3396), .IN5(n1827), 
        .Q(n1824) );
  OA22X1 U923 ( .IN1(n30), .IN2(n3393), .IN3(n990), .IN4(n3390), .Q(n1827) );
  OA221X1 U924 ( .IN1(n798), .IN2(n3387), .IN3(n830), .IN4(n3384), .IN5(n1828), 
        .Q(n1823) );
  OA22X1 U925 ( .IN1(n894), .IN2(n3381), .IN3(n862), .IN4(n3378), .Q(n1828) );
  OA221X1 U926 ( .IN1(n734), .IN2(n3375), .IN3(n766), .IN4(n3372), .IN5(n1829), 
        .Q(n1822) );
  OA22X1 U927 ( .IN1(n702), .IN2(n3369), .IN3(n670), .IN4(n3366), .Q(n1829) );
  OR2X1 U928 ( .IN1(n1830), .IN2(n1831), .Q(rd_dataA[29]) );
  NAND4X0 U929 ( .IN1(n1832), .IN2(n1833), .IN3(n1834), .IN4(n1835), .QN(n1831) );
  OA221X1 U930 ( .IN1(n515), .IN2(n3456), .IN3(n547), .IN4(n3453), .IN5(n1836), 
        .Q(n1835) );
  OA22X1 U931 ( .IN1(n611), .IN2(n3450), .IN3(n579), .IN4(n3447), .Q(n1836) );
  OA221X1 U932 ( .IN1(n387), .IN2(n3444), .IN3(n419), .IN4(n3441), .IN5(n1837), 
        .Q(n1834) );
  OA22X1 U933 ( .IN1(n483), .IN2(n3438), .IN3(n451), .IN4(n3435), .Q(n1837) );
  OA221X1 U934 ( .IN1(n259), .IN2(n3432), .IN3(n291), .IN4(n3429), .IN5(n1838), 
        .Q(n1833) );
  OA22X1 U935 ( .IN1(n355), .IN2(n3426), .IN3(n323), .IN4(n3423), .Q(n1838) );
  OA222X1 U936 ( .IN1(n163), .IN2(n3420), .IN3(n227), .IN4(n3417), .IN5(n195), 
        .IN6(n3414), .Q(n1832) );
  NAND4X0 U937 ( .IN1(n1839), .IN2(n1840), .IN3(n1841), .IN4(n1842), .QN(n1830) );
  OA221X1 U938 ( .IN1(n99), .IN2(n3411), .IN3(n67), .IN4(n3408), .IN5(n1843), 
        .Q(n1842) );
  OA22X1 U939 ( .IN1(n131), .IN2(n3405), .IN3(n35), .IN4(n3402), .Q(n1843) );
  OA221X1 U940 ( .IN1(n899), .IN2(n3399), .IN3(n931), .IN4(n3396), .IN5(n1844), 
        .Q(n1841) );
  OA22X1 U941 ( .IN1(n3), .IN2(n3393), .IN3(n963), .IN4(n3390), .Q(n1844) );
  OA221X1 U942 ( .IN1(n771), .IN2(n3387), .IN3(n803), .IN4(n3384), .IN5(n1845), 
        .Q(n1840) );
  OA22X1 U943 ( .IN1(n867), .IN2(n3381), .IN3(n835), .IN4(n3378), .Q(n1845) );
  OA221X1 U944 ( .IN1(n707), .IN2(n3375), .IN3(n739), .IN4(n3372), .IN5(n1846), 
        .Q(n1839) );
  OA22X1 U945 ( .IN1(n675), .IN2(n3369), .IN3(n643), .IN4(n3366), .Q(n1846) );
  OR2X1 U946 ( .IN1(n1847), .IN2(n1848), .Q(rd_dataA[28]) );
  NAND4X0 U947 ( .IN1(n1849), .IN2(n1850), .IN3(n1851), .IN4(n1852), .QN(n1848) );
  OA221X1 U948 ( .IN1(n516), .IN2(n3456), .IN3(n548), .IN4(n3453), .IN5(n1853), 
        .Q(n1852) );
  OA22X1 U949 ( .IN1(n612), .IN2(n3450), .IN3(n580), .IN4(n3447), .Q(n1853) );
  OA221X1 U950 ( .IN1(n388), .IN2(n3444), .IN3(n420), .IN4(n3441), .IN5(n1854), 
        .Q(n1851) );
  OA22X1 U951 ( .IN1(n484), .IN2(n3438), .IN3(n452), .IN4(n3435), .Q(n1854) );
  OA221X1 U952 ( .IN1(n260), .IN2(n3432), .IN3(n292), .IN4(n3429), .IN5(n1855), 
        .Q(n1850) );
  OA22X1 U953 ( .IN1(n356), .IN2(n3426), .IN3(n324), .IN4(n3423), .Q(n1855) );
  OA222X1 U954 ( .IN1(n164), .IN2(n3420), .IN3(n228), .IN4(n3417), .IN5(n196), 
        .IN6(n3414), .Q(n1849) );
  NAND4X0 U955 ( .IN1(n1856), .IN2(n1857), .IN3(n1858), .IN4(n1859), .QN(n1847) );
  OA221X1 U956 ( .IN1(n100), .IN2(n3411), .IN3(n68), .IN4(n3408), .IN5(n1860), 
        .Q(n1859) );
  OA22X1 U957 ( .IN1(n132), .IN2(n3405), .IN3(n36), .IN4(n3402), .Q(n1860) );
  OA221X1 U958 ( .IN1(n900), .IN2(n3399), .IN3(n932), .IN4(n3396), .IN5(n1861), 
        .Q(n1858) );
  OA22X1 U959 ( .IN1(n4), .IN2(n3393), .IN3(n964), .IN4(n3390), .Q(n1861) );
  OA221X1 U960 ( .IN1(n772), .IN2(n3387), .IN3(n804), .IN4(n3384), .IN5(n1862), 
        .Q(n1857) );
  OA22X1 U961 ( .IN1(n868), .IN2(n3381), .IN3(n836), .IN4(n3378), .Q(n1862) );
  OA221X1 U962 ( .IN1(n708), .IN2(n3375), .IN3(n740), .IN4(n3372), .IN5(n1863), 
        .Q(n1856) );
  OA22X1 U963 ( .IN1(n676), .IN2(n3369), .IN3(n644), .IN4(n3366), .Q(n1863) );
  OR2X1 U964 ( .IN1(n1864), .IN2(n1865), .Q(rd_dataA[27]) );
  NAND4X0 U965 ( .IN1(n1866), .IN2(n1867), .IN3(n1868), .IN4(n1869), .QN(n1865) );
  OA221X1 U966 ( .IN1(n517), .IN2(n3457), .IN3(n549), .IN4(n3454), .IN5(n1870), 
        .Q(n1869) );
  OA22X1 U967 ( .IN1(n613), .IN2(n3451), .IN3(n581), .IN4(n3448), .Q(n1870) );
  OA221X1 U968 ( .IN1(n389), .IN2(n3445), .IN3(n421), .IN4(n3442), .IN5(n1871), 
        .Q(n1868) );
  OA22X1 U969 ( .IN1(n485), .IN2(n3439), .IN3(n453), .IN4(n3436), .Q(n1871) );
  OA221X1 U970 ( .IN1(n261), .IN2(n3433), .IN3(n293), .IN4(n3430), .IN5(n1872), 
        .Q(n1867) );
  OA22X1 U971 ( .IN1(n357), .IN2(n3427), .IN3(n325), .IN4(n3424), .Q(n1872) );
  OA222X1 U972 ( .IN1(n165), .IN2(n3421), .IN3(n229), .IN4(n3418), .IN5(n197), 
        .IN6(n3415), .Q(n1866) );
  NAND4X0 U973 ( .IN1(n1873), .IN2(n1874), .IN3(n1875), .IN4(n1876), .QN(n1864) );
  OA221X1 U974 ( .IN1(n101), .IN2(n3412), .IN3(n69), .IN4(n3409), .IN5(n1877), 
        .Q(n1876) );
  OA22X1 U975 ( .IN1(n133), .IN2(n3406), .IN3(n37), .IN4(n3403), .Q(n1877) );
  OA221X1 U976 ( .IN1(n901), .IN2(n3400), .IN3(n933), .IN4(n3397), .IN5(n1878), 
        .Q(n1875) );
  OA22X1 U977 ( .IN1(n5), .IN2(n3394), .IN3(n965), .IN4(n3391), .Q(n1878) );
  OA221X1 U978 ( .IN1(n773), .IN2(n3388), .IN3(n805), .IN4(n3385), .IN5(n1879), 
        .Q(n1874) );
  OA22X1 U979 ( .IN1(n869), .IN2(n3382), .IN3(n837), .IN4(n3379), .Q(n1879) );
  OA221X1 U980 ( .IN1(n709), .IN2(n3376), .IN3(n741), .IN4(n3373), .IN5(n1880), 
        .Q(n1873) );
  OA22X1 U981 ( .IN1(n677), .IN2(n3370), .IN3(n645), .IN4(n3367), .Q(n1880) );
  OR2X1 U982 ( .IN1(n1881), .IN2(n1882), .Q(rd_dataA[26]) );
  NAND4X0 U983 ( .IN1(n1883), .IN2(n1884), .IN3(n1885), .IN4(n1886), .QN(n1882) );
  OA221X1 U984 ( .IN1(n518), .IN2(n3457), .IN3(n550), .IN4(n3454), .IN5(n1887), 
        .Q(n1886) );
  OA22X1 U985 ( .IN1(n614), .IN2(n3451), .IN3(n582), .IN4(n3448), .Q(n1887) );
  OA221X1 U986 ( .IN1(n390), .IN2(n3445), .IN3(n422), .IN4(n3442), .IN5(n1888), 
        .Q(n1885) );
  OA22X1 U987 ( .IN1(n486), .IN2(n3439), .IN3(n454), .IN4(n3436), .Q(n1888) );
  OA221X1 U988 ( .IN1(n262), .IN2(n3433), .IN3(n294), .IN4(n3430), .IN5(n1889), 
        .Q(n1884) );
  OA22X1 U989 ( .IN1(n358), .IN2(n3427), .IN3(n326), .IN4(n3424), .Q(n1889) );
  OA222X1 U990 ( .IN1(n166), .IN2(n3421), .IN3(n230), .IN4(n3418), .IN5(n198), 
        .IN6(n3415), .Q(n1883) );
  NAND4X0 U991 ( .IN1(n1890), .IN2(n1891), .IN3(n1892), .IN4(n1893), .QN(n1881) );
  OA221X1 U992 ( .IN1(n102), .IN2(n3412), .IN3(n70), .IN4(n3409), .IN5(n1894), 
        .Q(n1893) );
  OA22X1 U993 ( .IN1(n134), .IN2(n3406), .IN3(n38), .IN4(n3403), .Q(n1894) );
  OA221X1 U994 ( .IN1(n902), .IN2(n3400), .IN3(n934), .IN4(n3397), .IN5(n1895), 
        .Q(n1892) );
  OA22X1 U995 ( .IN1(n6), .IN2(n3394), .IN3(n966), .IN4(n3391), .Q(n1895) );
  OA221X1 U996 ( .IN1(n774), .IN2(n3388), .IN3(n806), .IN4(n3385), .IN5(n1896), 
        .Q(n1891) );
  OA22X1 U997 ( .IN1(n870), .IN2(n3382), .IN3(n838), .IN4(n3379), .Q(n1896) );
  OA221X1 U998 ( .IN1(n710), .IN2(n3376), .IN3(n742), .IN4(n3373), .IN5(n1897), 
        .Q(n1890) );
  OA22X1 U999 ( .IN1(n678), .IN2(n3370), .IN3(n646), .IN4(n3367), .Q(n1897) );
  OR2X1 U1000 ( .IN1(n1898), .IN2(n1899), .Q(rd_dataA[25]) );
  NAND4X0 U1001 ( .IN1(n1900), .IN2(n1901), .IN3(n1902), .IN4(n1903), .QN(
        n1899) );
  OA221X1 U1002 ( .IN1(n519), .IN2(n3457), .IN3(n551), .IN4(n3454), .IN5(n1904), .Q(n1903) );
  OA22X1 U1003 ( .IN1(n615), .IN2(n3451), .IN3(n583), .IN4(n3448), .Q(n1904)
         );
  OA221X1 U1004 ( .IN1(n391), .IN2(n3445), .IN3(n423), .IN4(n3442), .IN5(n1905), .Q(n1902) );
  OA22X1 U1005 ( .IN1(n487), .IN2(n3439), .IN3(n455), .IN4(n3436), .Q(n1905)
         );
  OA221X1 U1006 ( .IN1(n263), .IN2(n3433), .IN3(n295), .IN4(n3430), .IN5(n1906), .Q(n1901) );
  OA22X1 U1007 ( .IN1(n359), .IN2(n3427), .IN3(n327), .IN4(n3424), .Q(n1906)
         );
  OA222X1 U1008 ( .IN1(n167), .IN2(n3421), .IN3(n231), .IN4(n3418), .IN5(n199), 
        .IN6(n3415), .Q(n1900) );
  NAND4X0 U1009 ( .IN1(n1907), .IN2(n1908), .IN3(n1909), .IN4(n1910), .QN(
        n1898) );
  OA221X1 U1010 ( .IN1(n103), .IN2(n3412), .IN3(n71), .IN4(n3409), .IN5(n1911), 
        .Q(n1910) );
  OA22X1 U1011 ( .IN1(n135), .IN2(n3406), .IN3(n39), .IN4(n3403), .Q(n1911) );
  OA221X1 U1012 ( .IN1(n903), .IN2(n3400), .IN3(n935), .IN4(n3397), .IN5(n1912), .Q(n1909) );
  OA22X1 U1013 ( .IN1(n7), .IN2(n3394), .IN3(n967), .IN4(n3391), .Q(n1912) );
  OA221X1 U1014 ( .IN1(n775), .IN2(n3388), .IN3(n807), .IN4(n3385), .IN5(n1913), .Q(n1908) );
  OA22X1 U1015 ( .IN1(n871), .IN2(n3382), .IN3(n839), .IN4(n3379), .Q(n1913)
         );
  OA221X1 U1016 ( .IN1(n711), .IN2(n3376), .IN3(n743), .IN4(n3373), .IN5(n1914), .Q(n1907) );
  OA22X1 U1017 ( .IN1(n679), .IN2(n3370), .IN3(n647), .IN4(n3367), .Q(n1914)
         );
  OR2X1 U1018 ( .IN1(n1915), .IN2(n1916), .Q(rd_dataA[24]) );
  NAND4X0 U1019 ( .IN1(n1917), .IN2(n1918), .IN3(n1919), .IN4(n1920), .QN(
        n1916) );
  OA221X1 U1020 ( .IN1(n520), .IN2(n3457), .IN3(n552), .IN4(n3454), .IN5(n1921), .Q(n1920) );
  OA22X1 U1021 ( .IN1(n616), .IN2(n3451), .IN3(n584), .IN4(n3448), .Q(n1921)
         );
  OA221X1 U1022 ( .IN1(n392), .IN2(n3445), .IN3(n424), .IN4(n3442), .IN5(n1922), .Q(n1919) );
  OA22X1 U1023 ( .IN1(n488), .IN2(n3439), .IN3(n456), .IN4(n3436), .Q(n1922)
         );
  OA221X1 U1024 ( .IN1(n264), .IN2(n3433), .IN3(n296), .IN4(n3430), .IN5(n1923), .Q(n1918) );
  OA22X1 U1025 ( .IN1(n360), .IN2(n3427), .IN3(n328), .IN4(n3424), .Q(n1923)
         );
  OA222X1 U1026 ( .IN1(n168), .IN2(n3421), .IN3(n232), .IN4(n3418), .IN5(n200), 
        .IN6(n3415), .Q(n1917) );
  NAND4X0 U1027 ( .IN1(n1924), .IN2(n1925), .IN3(n1926), .IN4(n1927), .QN(
        n1915) );
  OA221X1 U1028 ( .IN1(n104), .IN2(n3412), .IN3(n72), .IN4(n3409), .IN5(n1928), 
        .Q(n1927) );
  OA22X1 U1029 ( .IN1(n136), .IN2(n3406), .IN3(n40), .IN4(n3403), .Q(n1928) );
  OA221X1 U1030 ( .IN1(n904), .IN2(n3400), .IN3(n936), .IN4(n3397), .IN5(n1929), .Q(n1926) );
  OA22X1 U1031 ( .IN1(n8), .IN2(n3394), .IN3(n968), .IN4(n3391), .Q(n1929) );
  OA221X1 U1032 ( .IN1(n776), .IN2(n3388), .IN3(n808), .IN4(n3385), .IN5(n1930), .Q(n1925) );
  OA22X1 U1033 ( .IN1(n872), .IN2(n3382), .IN3(n840), .IN4(n3379), .Q(n1930)
         );
  OA221X1 U1034 ( .IN1(n712), .IN2(n3376), .IN3(n744), .IN4(n3373), .IN5(n1931), .Q(n1924) );
  OA22X1 U1035 ( .IN1(n680), .IN2(n3370), .IN3(n648), .IN4(n3367), .Q(n1931)
         );
  OR2X1 U1036 ( .IN1(n1932), .IN2(n1933), .Q(rd_dataA[23]) );
  NAND4X0 U1037 ( .IN1(n1934), .IN2(n1935), .IN3(n1936), .IN4(n1937), .QN(
        n1933) );
  OA221X1 U1038 ( .IN1(n521), .IN2(n3457), .IN3(n553), .IN4(n3454), .IN5(n1938), .Q(n1937) );
  OA22X1 U1039 ( .IN1(n617), .IN2(n3451), .IN3(n585), .IN4(n3448), .Q(n1938)
         );
  OA221X1 U1040 ( .IN1(n393), .IN2(n3445), .IN3(n425), .IN4(n3442), .IN5(n1939), .Q(n1936) );
  OA22X1 U1041 ( .IN1(n489), .IN2(n3439), .IN3(n457), .IN4(n3436), .Q(n1939)
         );
  OA221X1 U1042 ( .IN1(n265), .IN2(n3433), .IN3(n297), .IN4(n3430), .IN5(n1940), .Q(n1935) );
  OA22X1 U1043 ( .IN1(n361), .IN2(n3427), .IN3(n329), .IN4(n3424), .Q(n1940)
         );
  OA222X1 U1044 ( .IN1(n169), .IN2(n3421), .IN3(n233), .IN4(n3418), .IN5(n201), 
        .IN6(n3415), .Q(n1934) );
  NAND4X0 U1045 ( .IN1(n1941), .IN2(n1942), .IN3(n1943), .IN4(n1944), .QN(
        n1932) );
  OA221X1 U1046 ( .IN1(n105), .IN2(n3412), .IN3(n73), .IN4(n3409), .IN5(n1945), 
        .Q(n1944) );
  OA22X1 U1047 ( .IN1(n137), .IN2(n3406), .IN3(n41), .IN4(n3403), .Q(n1945) );
  OA221X1 U1048 ( .IN1(n905), .IN2(n3400), .IN3(n937), .IN4(n3397), .IN5(n1946), .Q(n1943) );
  OA22X1 U1049 ( .IN1(n9), .IN2(n3394), .IN3(n969), .IN4(n3391), .Q(n1946) );
  OA221X1 U1050 ( .IN1(n777), .IN2(n3388), .IN3(n809), .IN4(n3385), .IN5(n1947), .Q(n1942) );
  OA22X1 U1051 ( .IN1(n873), .IN2(n3382), .IN3(n841), .IN4(n3379), .Q(n1947)
         );
  OA221X1 U1052 ( .IN1(n713), .IN2(n3376), .IN3(n745), .IN4(n3373), .IN5(n1948), .Q(n1941) );
  OA22X1 U1053 ( .IN1(n681), .IN2(n3370), .IN3(n649), .IN4(n3367), .Q(n1948)
         );
  OR2X1 U1054 ( .IN1(n1949), .IN2(n1950), .Q(rd_dataA[22]) );
  NAND4X0 U1055 ( .IN1(n1951), .IN2(n1952), .IN3(n1953), .IN4(n1954), .QN(
        n1950) );
  OA221X1 U1056 ( .IN1(n522), .IN2(n3457), .IN3(n554), .IN4(n3454), .IN5(n1955), .Q(n1954) );
  OA22X1 U1057 ( .IN1(n618), .IN2(n3451), .IN3(n586), .IN4(n3448), .Q(n1955)
         );
  OA221X1 U1058 ( .IN1(n394), .IN2(n3445), .IN3(n426), .IN4(n3442), .IN5(n1956), .Q(n1953) );
  OA22X1 U1059 ( .IN1(n490), .IN2(n3439), .IN3(n458), .IN4(n3436), .Q(n1956)
         );
  OA221X1 U1060 ( .IN1(n266), .IN2(n3433), .IN3(n298), .IN4(n3430), .IN5(n1957), .Q(n1952) );
  OA22X1 U1061 ( .IN1(n362), .IN2(n3427), .IN3(n330), .IN4(n3424), .Q(n1957)
         );
  OA222X1 U1062 ( .IN1(n170), .IN2(n3421), .IN3(n234), .IN4(n3418), .IN5(n202), 
        .IN6(n3415), .Q(n1951) );
  NAND4X0 U1063 ( .IN1(n1958), .IN2(n1959), .IN3(n1960), .IN4(n1961), .QN(
        n1949) );
  OA221X1 U1064 ( .IN1(n106), .IN2(n3412), .IN3(n74), .IN4(n3409), .IN5(n1962), 
        .Q(n1961) );
  OA22X1 U1065 ( .IN1(n138), .IN2(n3406), .IN3(n42), .IN4(n3403), .Q(n1962) );
  OA221X1 U1066 ( .IN1(n906), .IN2(n3400), .IN3(n938), .IN4(n3397), .IN5(n1963), .Q(n1960) );
  OA22X1 U1067 ( .IN1(n10), .IN2(n3394), .IN3(n970), .IN4(n3391), .Q(n1963) );
  OA221X1 U1068 ( .IN1(n778), .IN2(n3388), .IN3(n810), .IN4(n3385), .IN5(n1964), .Q(n1959) );
  OA22X1 U1069 ( .IN1(n874), .IN2(n3382), .IN3(n842), .IN4(n3379), .Q(n1964)
         );
  OA221X1 U1070 ( .IN1(n714), .IN2(n3376), .IN3(n746), .IN4(n3373), .IN5(n1965), .Q(n1958) );
  OA22X1 U1071 ( .IN1(n682), .IN2(n3370), .IN3(n650), .IN4(n3367), .Q(n1965)
         );
  OR2X1 U1072 ( .IN1(n1966), .IN2(n1967), .Q(rd_dataA[21]) );
  NAND4X0 U1073 ( .IN1(n1968), .IN2(n1969), .IN3(n1970), .IN4(n1971), .QN(
        n1967) );
  OA221X1 U1074 ( .IN1(n523), .IN2(n3457), .IN3(n555), .IN4(n3454), .IN5(n1972), .Q(n1971) );
  OA22X1 U1075 ( .IN1(n619), .IN2(n3451), .IN3(n587), .IN4(n3448), .Q(n1972)
         );
  OA221X1 U1076 ( .IN1(n395), .IN2(n3445), .IN3(n427), .IN4(n3442), .IN5(n1973), .Q(n1970) );
  OA22X1 U1077 ( .IN1(n491), .IN2(n3439), .IN3(n459), .IN4(n3436), .Q(n1973)
         );
  OA221X1 U1078 ( .IN1(n267), .IN2(n3433), .IN3(n299), .IN4(n3430), .IN5(n1974), .Q(n1969) );
  OA22X1 U1079 ( .IN1(n363), .IN2(n3427), .IN3(n331), .IN4(n3424), .Q(n1974)
         );
  OA222X1 U1080 ( .IN1(n171), .IN2(n3421), .IN3(n235), .IN4(n3418), .IN5(n203), 
        .IN6(n3415), .Q(n1968) );
  NAND4X0 U1081 ( .IN1(n1975), .IN2(n1976), .IN3(n1977), .IN4(n1978), .QN(
        n1966) );
  OA221X1 U1082 ( .IN1(n107), .IN2(n3412), .IN3(n75), .IN4(n3409), .IN5(n1979), 
        .Q(n1978) );
  OA22X1 U1083 ( .IN1(n139), .IN2(n3406), .IN3(n43), .IN4(n3403), .Q(n1979) );
  OA221X1 U1084 ( .IN1(n907), .IN2(n3400), .IN3(n939), .IN4(n3397), .IN5(n1980), .Q(n1977) );
  OA22X1 U1085 ( .IN1(n11), .IN2(n3394), .IN3(n971), .IN4(n3391), .Q(n1980) );
  OA221X1 U1086 ( .IN1(n779), .IN2(n3388), .IN3(n811), .IN4(n3385), .IN5(n1981), .Q(n1976) );
  OA22X1 U1087 ( .IN1(n875), .IN2(n3382), .IN3(n843), .IN4(n3379), .Q(n1981)
         );
  OA221X1 U1088 ( .IN1(n715), .IN2(n3376), .IN3(n747), .IN4(n3373), .IN5(n1982), .Q(n1975) );
  OA22X1 U1089 ( .IN1(n683), .IN2(n3370), .IN3(n651), .IN4(n3367), .Q(n1982)
         );
  OR2X1 U1090 ( .IN1(n1983), .IN2(n1984), .Q(rd_dataA[20]) );
  NAND4X0 U1091 ( .IN1(n1985), .IN2(n1986), .IN3(n1987), .IN4(n1988), .QN(
        n1984) );
  OA221X1 U1092 ( .IN1(n524), .IN2(n3457), .IN3(n556), .IN4(n3454), .IN5(n1989), .Q(n1988) );
  OA22X1 U1093 ( .IN1(n620), .IN2(n3451), .IN3(n588), .IN4(n3448), .Q(n1989)
         );
  OA221X1 U1094 ( .IN1(n396), .IN2(n3445), .IN3(n428), .IN4(n3442), .IN5(n1990), .Q(n1987) );
  OA22X1 U1095 ( .IN1(n492), .IN2(n3439), .IN3(n460), .IN4(n3436), .Q(n1990)
         );
  OA221X1 U1096 ( .IN1(n268), .IN2(n3433), .IN3(n300), .IN4(n3430), .IN5(n1991), .Q(n1986) );
  OA22X1 U1097 ( .IN1(n364), .IN2(n3427), .IN3(n332), .IN4(n3424), .Q(n1991)
         );
  OA222X1 U1098 ( .IN1(n172), .IN2(n3421), .IN3(n236), .IN4(n3418), .IN5(n204), 
        .IN6(n3415), .Q(n1985) );
  NAND4X0 U1099 ( .IN1(n1992), .IN2(n1993), .IN3(n1994), .IN4(n1995), .QN(
        n1983) );
  OA221X1 U1100 ( .IN1(n108), .IN2(n3412), .IN3(n76), .IN4(n3409), .IN5(n1996), 
        .Q(n1995) );
  OA22X1 U1101 ( .IN1(n140), .IN2(n3406), .IN3(n44), .IN4(n3403), .Q(n1996) );
  OA221X1 U1102 ( .IN1(n908), .IN2(n3400), .IN3(n940), .IN4(n3397), .IN5(n1997), .Q(n1994) );
  OA22X1 U1103 ( .IN1(n12), .IN2(n3394), .IN3(n972), .IN4(n3391), .Q(n1997) );
  OA221X1 U1104 ( .IN1(n780), .IN2(n3388), .IN3(n812), .IN4(n3385), .IN5(n1998), .Q(n1993) );
  OA22X1 U1105 ( .IN1(n876), .IN2(n3382), .IN3(n844), .IN4(n3379), .Q(n1998)
         );
  OA221X1 U1106 ( .IN1(n716), .IN2(n3376), .IN3(n748), .IN4(n3373), .IN5(n1999), .Q(n1992) );
  OA22X1 U1107 ( .IN1(n684), .IN2(n3370), .IN3(n652), .IN4(n3367), .Q(n1999)
         );
  OA221X1 U1110 ( .IN1(n543), .IN2(n3457), .IN3(n575), .IN4(n3454), .IN5(n2006), .Q(n2005) );
  OA22X1 U1111 ( .IN1(n639), .IN2(n3451), .IN3(n607), .IN4(n3448), .Q(n2006)
         );
  OA221X1 U1112 ( .IN1(n415), .IN2(n3445), .IN3(n447), .IN4(n3442), .IN5(n2007), .Q(n2004) );
  OA22X1 U1113 ( .IN1(n511), .IN2(n3439), .IN3(n479), .IN4(n3436), .Q(n2007)
         );
  OA221X1 U1114 ( .IN1(n287), .IN2(n3433), .IN3(n319), .IN4(n3430), .IN5(n2008), .Q(n2003) );
  OA22X1 U1115 ( .IN1(n383), .IN2(n3427), .IN3(n351), .IN4(n3424), .Q(n2008)
         );
  OA222X1 U1116 ( .IN1(n191), .IN2(n3421), .IN3(n255), .IN4(n3418), .IN5(n223), 
        .IN6(n3415), .Q(n2002) );
  OA221X1 U1118 ( .IN1(n127), .IN2(n3412), .IN3(n95), .IN4(n3409), .IN5(n2013), 
        .Q(n2012) );
  OA22X1 U1119 ( .IN1(n159), .IN2(n3406), .IN3(n63), .IN4(n3403), .Q(n2013) );
  OA221X1 U1120 ( .IN1(n927), .IN2(n3400), .IN3(n959), .IN4(n3397), .IN5(n2014), .Q(n2011) );
  OA22X1 U1121 ( .IN1(n31), .IN2(n3394), .IN3(n991), .IN4(n3391), .Q(n2014) );
  OA221X1 U1122 ( .IN1(n799), .IN2(n3388), .IN3(n831), .IN4(n3385), .IN5(n2015), .Q(n2010) );
  OA22X1 U1123 ( .IN1(n895), .IN2(n3382), .IN3(n863), .IN4(n3379), .Q(n2015)
         );
  OA221X1 U1124 ( .IN1(n735), .IN2(n3376), .IN3(n767), .IN4(n3373), .IN5(n2016), .Q(n2009) );
  OA22X1 U1125 ( .IN1(n703), .IN2(n3370), .IN3(n671), .IN4(n3367), .Q(n2016)
         );
  OR2X1 U1126 ( .IN1(n2017), .IN2(n2018), .Q(rd_dataA[19]) );
  NAND4X0 U1127 ( .IN1(n2019), .IN2(n2020), .IN3(n2021), .IN4(n2022), .QN(
        n2018) );
  OA221X1 U1128 ( .IN1(n525), .IN2(n3457), .IN3(n557), .IN4(n3454), .IN5(n2023), .Q(n2022) );
  OA22X1 U1129 ( .IN1(n621), .IN2(n3451), .IN3(n589), .IN4(n3448), .Q(n2023)
         );
  OA221X1 U1130 ( .IN1(n397), .IN2(n3445), .IN3(n429), .IN4(n3442), .IN5(n2024), .Q(n2021) );
  OA22X1 U1131 ( .IN1(n493), .IN2(n3439), .IN3(n461), .IN4(n3436), .Q(n2024)
         );
  OA221X1 U1132 ( .IN1(n269), .IN2(n3433), .IN3(n301), .IN4(n3430), .IN5(n2025), .Q(n2020) );
  OA22X1 U1133 ( .IN1(n365), .IN2(n3427), .IN3(n333), .IN4(n3424), .Q(n2025)
         );
  OA222X1 U1134 ( .IN1(n173), .IN2(n3421), .IN3(n237), .IN4(n3418), .IN5(n205), 
        .IN6(n3415), .Q(n2019) );
  NAND4X0 U1135 ( .IN1(n2026), .IN2(n2027), .IN3(n2028), .IN4(n2029), .QN(
        n2017) );
  OA221X1 U1136 ( .IN1(n109), .IN2(n3412), .IN3(n77), .IN4(n3409), .IN5(n2030), 
        .Q(n2029) );
  OA22X1 U1137 ( .IN1(n141), .IN2(n3406), .IN3(n45), .IN4(n3403), .Q(n2030) );
  OA221X1 U1138 ( .IN1(n909), .IN2(n3400), .IN3(n941), .IN4(n3397), .IN5(n2031), .Q(n2028) );
  OA22X1 U1139 ( .IN1(n13), .IN2(n3394), .IN3(n973), .IN4(n3391), .Q(n2031) );
  OA221X1 U1140 ( .IN1(n781), .IN2(n3388), .IN3(n813), .IN4(n3385), .IN5(n2032), .Q(n2027) );
  OA22X1 U1141 ( .IN1(n877), .IN2(n3382), .IN3(n845), .IN4(n3379), .Q(n2032)
         );
  OA221X1 U1142 ( .IN1(n717), .IN2(n3376), .IN3(n749), .IN4(n3373), .IN5(n2033), .Q(n2026) );
  OA22X1 U1143 ( .IN1(n685), .IN2(n3370), .IN3(n653), .IN4(n3367), .Q(n2033)
         );
  OR2X1 U1144 ( .IN1(n2034), .IN2(n2035), .Q(rd_dataA[18]) );
  NAND4X0 U1145 ( .IN1(n2036), .IN2(n2037), .IN3(n2038), .IN4(n2039), .QN(
        n2035) );
  OA221X1 U1146 ( .IN1(n526), .IN2(n3457), .IN3(n558), .IN4(n3454), .IN5(n2040), .Q(n2039) );
  OA22X1 U1147 ( .IN1(n622), .IN2(n3451), .IN3(n590), .IN4(n3448), .Q(n2040)
         );
  OA221X1 U1148 ( .IN1(n398), .IN2(n3445), .IN3(n430), .IN4(n3442), .IN5(n2041), .Q(n2038) );
  OA22X1 U1149 ( .IN1(n494), .IN2(n3439), .IN3(n462), .IN4(n3436), .Q(n2041)
         );
  OA221X1 U1150 ( .IN1(n270), .IN2(n3433), .IN3(n302), .IN4(n3430), .IN5(n2042), .Q(n2037) );
  OA22X1 U1151 ( .IN1(n366), .IN2(n3427), .IN3(n334), .IN4(n3424), .Q(n2042)
         );
  OA222X1 U1152 ( .IN1(n174), .IN2(n3421), .IN3(n238), .IN4(n3418), .IN5(n206), 
        .IN6(n3415), .Q(n2036) );
  NAND4X0 U1153 ( .IN1(n2043), .IN2(n2044), .IN3(n2045), .IN4(n2046), .QN(
        n2034) );
  OA221X1 U1154 ( .IN1(n110), .IN2(n3412), .IN3(n78), .IN4(n3409), .IN5(n2047), 
        .Q(n2046) );
  OA22X1 U1155 ( .IN1(n142), .IN2(n3406), .IN3(n46), .IN4(n3403), .Q(n2047) );
  OA221X1 U1156 ( .IN1(n910), .IN2(n3400), .IN3(n942), .IN4(n3397), .IN5(n2048), .Q(n2045) );
  OA22X1 U1157 ( .IN1(n14), .IN2(n3394), .IN3(n974), .IN4(n3391), .Q(n2048) );
  OA221X1 U1158 ( .IN1(n782), .IN2(n3388), .IN3(n814), .IN4(n3385), .IN5(n2049), .Q(n2044) );
  OA22X1 U1159 ( .IN1(n878), .IN2(n3382), .IN3(n846), .IN4(n3379), .Q(n2049)
         );
  OA221X1 U1160 ( .IN1(n718), .IN2(n3376), .IN3(n750), .IN4(n3373), .IN5(n2050), .Q(n2043) );
  OA22X1 U1161 ( .IN1(n686), .IN2(n3370), .IN3(n654), .IN4(n3367), .Q(n2050)
         );
  OR2X1 U1162 ( .IN1(n2051), .IN2(n2052), .Q(rd_dataA[17]) );
  NAND4X0 U1163 ( .IN1(n2053), .IN2(n2054), .IN3(n2055), .IN4(n2056), .QN(
        n2052) );
  OA221X1 U1164 ( .IN1(n527), .IN2(n3457), .IN3(n559), .IN4(n3454), .IN5(n2057), .Q(n2056) );
  OA22X1 U1165 ( .IN1(n623), .IN2(n3451), .IN3(n591), .IN4(n3448), .Q(n2057)
         );
  OA221X1 U1166 ( .IN1(n399), .IN2(n3445), .IN3(n431), .IN4(n3442), .IN5(n2058), .Q(n2055) );
  OA22X1 U1167 ( .IN1(n495), .IN2(n3439), .IN3(n463), .IN4(n3436), .Q(n2058)
         );
  OA221X1 U1168 ( .IN1(n271), .IN2(n3433), .IN3(n303), .IN4(n3430), .IN5(n2059), .Q(n2054) );
  OA22X1 U1169 ( .IN1(n367), .IN2(n3427), .IN3(n335), .IN4(n3424), .Q(n2059)
         );
  OA222X1 U1170 ( .IN1(n175), .IN2(n3421), .IN3(n239), .IN4(n3418), .IN5(n207), 
        .IN6(n3415), .Q(n2053) );
  NAND4X0 U1171 ( .IN1(n2060), .IN2(n2061), .IN3(n2062), .IN4(n2063), .QN(
        n2051) );
  OA221X1 U1172 ( .IN1(n111), .IN2(n3412), .IN3(n79), .IN4(n3409), .IN5(n2064), 
        .Q(n2063) );
  OA22X1 U1173 ( .IN1(n143), .IN2(n3406), .IN3(n47), .IN4(n3403), .Q(n2064) );
  OA221X1 U1174 ( .IN1(n911), .IN2(n3400), .IN3(n943), .IN4(n3397), .IN5(n2065), .Q(n2062) );
  OA22X1 U1175 ( .IN1(n15), .IN2(n3394), .IN3(n975), .IN4(n3391), .Q(n2065) );
  OA221X1 U1176 ( .IN1(n783), .IN2(n3388), .IN3(n815), .IN4(n3385), .IN5(n2066), .Q(n2061) );
  OA22X1 U1177 ( .IN1(n879), .IN2(n3382), .IN3(n847), .IN4(n3379), .Q(n2066)
         );
  OA221X1 U1178 ( .IN1(n719), .IN2(n3376), .IN3(n751), .IN4(n3373), .IN5(n2067), .Q(n2060) );
  OA22X1 U1179 ( .IN1(n687), .IN2(n3370), .IN3(n655), .IN4(n3367), .Q(n2067)
         );
  OR2X1 U1180 ( .IN1(n2068), .IN2(n2069), .Q(rd_dataA[16]) );
  NAND4X0 U1181 ( .IN1(n2070), .IN2(n2071), .IN3(n2072), .IN4(n2073), .QN(
        n2069) );
  OA221X1 U1182 ( .IN1(n528), .IN2(n3458), .IN3(n560), .IN4(n3455), .IN5(n2074), .Q(n2073) );
  OA22X1 U1183 ( .IN1(n624), .IN2(n3452), .IN3(n592), .IN4(n3449), .Q(n2074)
         );
  OA221X1 U1184 ( .IN1(n400), .IN2(n3446), .IN3(n432), .IN4(n3443), .IN5(n2075), .Q(n2072) );
  OA22X1 U1185 ( .IN1(n496), .IN2(n3440), .IN3(n464), .IN4(n3437), .Q(n2075)
         );
  OA221X1 U1186 ( .IN1(n272), .IN2(n3434), .IN3(n304), .IN4(n3431), .IN5(n2076), .Q(n2071) );
  OA22X1 U1187 ( .IN1(n368), .IN2(n3428), .IN3(n336), .IN4(n3425), .Q(n2076)
         );
  OA222X1 U1188 ( .IN1(n176), .IN2(n3422), .IN3(n240), .IN4(n3419), .IN5(n208), 
        .IN6(n3416), .Q(n2070) );
  NAND4X0 U1189 ( .IN1(n2077), .IN2(n2078), .IN3(n2079), .IN4(n2080), .QN(
        n2068) );
  OA221X1 U1190 ( .IN1(n112), .IN2(n3413), .IN3(n80), .IN4(n3410), .IN5(n2081), 
        .Q(n2080) );
  OA22X1 U1191 ( .IN1(n144), .IN2(n3407), .IN3(n48), .IN4(n3404), .Q(n2081) );
  OA221X1 U1192 ( .IN1(n912), .IN2(n3401), .IN3(n944), .IN4(n3398), .IN5(n2082), .Q(n2079) );
  OA22X1 U1193 ( .IN1(n16), .IN2(n3395), .IN3(n976), .IN4(n3392), .Q(n2082) );
  OA221X1 U1194 ( .IN1(n784), .IN2(n3389), .IN3(n816), .IN4(n3386), .IN5(n2083), .Q(n2078) );
  OA22X1 U1195 ( .IN1(n880), .IN2(n3383), .IN3(n848), .IN4(n3380), .Q(n2083)
         );
  OA221X1 U1196 ( .IN1(n720), .IN2(n3377), .IN3(n752), .IN4(n3374), .IN5(n2084), .Q(n2077) );
  OA22X1 U1197 ( .IN1(n688), .IN2(n3371), .IN3(n656), .IN4(n3368), .Q(n2084)
         );
  OR2X1 U1198 ( .IN1(n2085), .IN2(n2086), .Q(rd_dataA[15]) );
  NAND4X0 U1199 ( .IN1(n2087), .IN2(n2088), .IN3(n2089), .IN4(n2090), .QN(
        n2086) );
  OA221X1 U1200 ( .IN1(n529), .IN2(n3458), .IN3(n561), .IN4(n3455), .IN5(n2091), .Q(n2090) );
  OA22X1 U1201 ( .IN1(n625), .IN2(n3452), .IN3(n593), .IN4(n3449), .Q(n2091)
         );
  OA221X1 U1202 ( .IN1(n401), .IN2(n3446), .IN3(n433), .IN4(n3443), .IN5(n2092), .Q(n2089) );
  OA22X1 U1203 ( .IN1(n497), .IN2(n3440), .IN3(n465), .IN4(n3437), .Q(n2092)
         );
  OA221X1 U1204 ( .IN1(n273), .IN2(n3434), .IN3(n305), .IN4(n3431), .IN5(n2093), .Q(n2088) );
  OA22X1 U1205 ( .IN1(n369), .IN2(n3428), .IN3(n337), .IN4(n3425), .Q(n2093)
         );
  OA222X1 U1206 ( .IN1(n177), .IN2(n3422), .IN3(n241), .IN4(n3419), .IN5(n209), 
        .IN6(n3416), .Q(n2087) );
  NAND4X0 U1207 ( .IN1(n2094), .IN2(n2095), .IN3(n2096), .IN4(n2097), .QN(
        n2085) );
  OA221X1 U1208 ( .IN1(n113), .IN2(n3413), .IN3(n81), .IN4(n3410), .IN5(n2098), 
        .Q(n2097) );
  OA22X1 U1209 ( .IN1(n145), .IN2(n3407), .IN3(n49), .IN4(n3404), .Q(n2098) );
  OA221X1 U1210 ( .IN1(n913), .IN2(n3401), .IN3(n945), .IN4(n3398), .IN5(n2099), .Q(n2096) );
  OA22X1 U1211 ( .IN1(n17), .IN2(n3395), .IN3(n977), .IN4(n3392), .Q(n2099) );
  OA221X1 U1212 ( .IN1(n785), .IN2(n3389), .IN3(n817), .IN4(n3386), .IN5(n2100), .Q(n2095) );
  OA22X1 U1213 ( .IN1(n881), .IN2(n3383), .IN3(n849), .IN4(n3380), .Q(n2100)
         );
  OA221X1 U1214 ( .IN1(n721), .IN2(n3377), .IN3(n753), .IN4(n3374), .IN5(n2101), .Q(n2094) );
  OA22X1 U1215 ( .IN1(n689), .IN2(n3371), .IN3(n657), .IN4(n3368), .Q(n2101)
         );
  OR2X1 U1216 ( .IN1(n2102), .IN2(n2103), .Q(rd_dataA[14]) );
  NAND4X0 U1217 ( .IN1(n2104), .IN2(n2105), .IN3(n2106), .IN4(n2107), .QN(
        n2103) );
  OA221X1 U1218 ( .IN1(n530), .IN2(n3458), .IN3(n562), .IN4(n3455), .IN5(n2108), .Q(n2107) );
  OA22X1 U1219 ( .IN1(n626), .IN2(n3452), .IN3(n594), .IN4(n3449), .Q(n2108)
         );
  OA221X1 U1220 ( .IN1(n402), .IN2(n3446), .IN3(n434), .IN4(n3443), .IN5(n2109), .Q(n2106) );
  OA22X1 U1221 ( .IN1(n498), .IN2(n3440), .IN3(n466), .IN4(n3437), .Q(n2109)
         );
  OA221X1 U1222 ( .IN1(n274), .IN2(n3434), .IN3(n306), .IN4(n3431), .IN5(n2110), .Q(n2105) );
  OA22X1 U1223 ( .IN1(n370), .IN2(n3428), .IN3(n338), .IN4(n3425), .Q(n2110)
         );
  OA222X1 U1224 ( .IN1(n178), .IN2(n3422), .IN3(n242), .IN4(n3419), .IN5(n210), 
        .IN6(n3416), .Q(n2104) );
  NAND4X0 U1225 ( .IN1(n2111), .IN2(n2112), .IN3(n2113), .IN4(n2114), .QN(
        n2102) );
  OA221X1 U1226 ( .IN1(n114), .IN2(n3413), .IN3(n82), .IN4(n3410), .IN5(n2115), 
        .Q(n2114) );
  OA22X1 U1227 ( .IN1(n146), .IN2(n3407), .IN3(n50), .IN4(n3404), .Q(n2115) );
  OA221X1 U1228 ( .IN1(n914), .IN2(n3401), .IN3(n946), .IN4(n3398), .IN5(n2116), .Q(n2113) );
  OA22X1 U1229 ( .IN1(n18), .IN2(n3395), .IN3(n978), .IN4(n3392), .Q(n2116) );
  OA221X1 U1230 ( .IN1(n786), .IN2(n3389), .IN3(n818), .IN4(n3386), .IN5(n2117), .Q(n2112) );
  OA22X1 U1231 ( .IN1(n882), .IN2(n3383), .IN3(n850), .IN4(n3380), .Q(n2117)
         );
  OA221X1 U1232 ( .IN1(n722), .IN2(n3377), .IN3(n754), .IN4(n3374), .IN5(n2118), .Q(n2111) );
  OA22X1 U1233 ( .IN1(n690), .IN2(n3371), .IN3(n658), .IN4(n3368), .Q(n2118)
         );
  OR2X1 U1234 ( .IN1(n2119), .IN2(n2120), .Q(rd_dataA[13]) );
  NAND4X0 U1235 ( .IN1(n2121), .IN2(n2122), .IN3(n2123), .IN4(n2124), .QN(
        n2120) );
  OA221X1 U1236 ( .IN1(n531), .IN2(n3458), .IN3(n563), .IN4(n3455), .IN5(n2125), .Q(n2124) );
  OA22X1 U1237 ( .IN1(n627), .IN2(n3452), .IN3(n595), .IN4(n3449), .Q(n2125)
         );
  OA221X1 U1238 ( .IN1(n403), .IN2(n3446), .IN3(n435), .IN4(n3443), .IN5(n2126), .Q(n2123) );
  OA22X1 U1239 ( .IN1(n499), .IN2(n3440), .IN3(n467), .IN4(n3437), .Q(n2126)
         );
  OA221X1 U1240 ( .IN1(n275), .IN2(n3434), .IN3(n307), .IN4(n3431), .IN5(n2127), .Q(n2122) );
  OA22X1 U1241 ( .IN1(n371), .IN2(n3428), .IN3(n339), .IN4(n3425), .Q(n2127)
         );
  OA222X1 U1242 ( .IN1(n179), .IN2(n3422), .IN3(n243), .IN4(n3419), .IN5(n211), 
        .IN6(n3416), .Q(n2121) );
  NAND4X0 U1243 ( .IN1(n2128), .IN2(n2129), .IN3(n2130), .IN4(n2131), .QN(
        n2119) );
  OA221X1 U1244 ( .IN1(n115), .IN2(n3413), .IN3(n83), .IN4(n3410), .IN5(n2132), 
        .Q(n2131) );
  OA22X1 U1245 ( .IN1(n147), .IN2(n3407), .IN3(n51), .IN4(n3404), .Q(n2132) );
  OA221X1 U1246 ( .IN1(n915), .IN2(n3401), .IN3(n947), .IN4(n3398), .IN5(n2133), .Q(n2130) );
  OA22X1 U1247 ( .IN1(n19), .IN2(n3395), .IN3(n979), .IN4(n3392), .Q(n2133) );
  OA221X1 U1248 ( .IN1(n787), .IN2(n3389), .IN3(n819), .IN4(n3386), .IN5(n2134), .Q(n2129) );
  OA22X1 U1249 ( .IN1(n883), .IN2(n3383), .IN3(n851), .IN4(n3380), .Q(n2134)
         );
  OA221X1 U1250 ( .IN1(n723), .IN2(n3377), .IN3(n755), .IN4(n3374), .IN5(n2135), .Q(n2128) );
  OA22X1 U1251 ( .IN1(n691), .IN2(n3371), .IN3(n659), .IN4(n3368), .Q(n2135)
         );
  OR2X1 U1252 ( .IN1(n2136), .IN2(n2137), .Q(rd_dataA[12]) );
  NAND4X0 U1253 ( .IN1(n2138), .IN2(n2139), .IN3(n2140), .IN4(n2141), .QN(
        n2137) );
  OA221X1 U1254 ( .IN1(n532), .IN2(n3458), .IN3(n564), .IN4(n3455), .IN5(n2142), .Q(n2141) );
  OA22X1 U1255 ( .IN1(n628), .IN2(n3452), .IN3(n596), .IN4(n3449), .Q(n2142)
         );
  OA221X1 U1256 ( .IN1(n404), .IN2(n3446), .IN3(n436), .IN4(n3443), .IN5(n2143), .Q(n2140) );
  OA22X1 U1257 ( .IN1(n500), .IN2(n3440), .IN3(n468), .IN4(n3437), .Q(n2143)
         );
  OA221X1 U1258 ( .IN1(n276), .IN2(n3434), .IN3(n308), .IN4(n3431), .IN5(n2144), .Q(n2139) );
  OA22X1 U1259 ( .IN1(n372), .IN2(n3428), .IN3(n340), .IN4(n3425), .Q(n2144)
         );
  OA222X1 U1260 ( .IN1(n180), .IN2(n3422), .IN3(n244), .IN4(n3419), .IN5(n212), 
        .IN6(n3416), .Q(n2138) );
  NAND4X0 U1261 ( .IN1(n2145), .IN2(n2146), .IN3(n2147), .IN4(n2148), .QN(
        n2136) );
  OA221X1 U1262 ( .IN1(n116), .IN2(n3413), .IN3(n84), .IN4(n3410), .IN5(n2149), 
        .Q(n2148) );
  OA22X1 U1263 ( .IN1(n148), .IN2(n3407), .IN3(n52), .IN4(n3404), .Q(n2149) );
  OA221X1 U1264 ( .IN1(n916), .IN2(n3401), .IN3(n948), .IN4(n3398), .IN5(n2150), .Q(n2147) );
  OA22X1 U1265 ( .IN1(n20), .IN2(n3395), .IN3(n980), .IN4(n3392), .Q(n2150) );
  OA221X1 U1266 ( .IN1(n788), .IN2(n3389), .IN3(n820), .IN4(n3386), .IN5(n2151), .Q(n2146) );
  OA22X1 U1267 ( .IN1(n884), .IN2(n3383), .IN3(n852), .IN4(n3380), .Q(n2151)
         );
  OA221X1 U1268 ( .IN1(n724), .IN2(n3377), .IN3(n756), .IN4(n3374), .IN5(n2152), .Q(n2145) );
  OA22X1 U1269 ( .IN1(n692), .IN2(n3371), .IN3(n660), .IN4(n3368), .Q(n2152)
         );
  OR2X1 U1270 ( .IN1(n2153), .IN2(n2154), .Q(rd_dataA[11]) );
  NAND4X0 U1271 ( .IN1(n2155), .IN2(n2156), .IN3(n2157), .IN4(n2158), .QN(
        n2154) );
  OA221X1 U1272 ( .IN1(n533), .IN2(n3458), .IN3(n565), .IN4(n3455), .IN5(n2159), .Q(n2158) );
  OA22X1 U1273 ( .IN1(n629), .IN2(n3452), .IN3(n597), .IN4(n3449), .Q(n2159)
         );
  OA221X1 U1274 ( .IN1(n405), .IN2(n3446), .IN3(n437), .IN4(n3443), .IN5(n2160), .Q(n2157) );
  OA22X1 U1275 ( .IN1(n501), .IN2(n3440), .IN3(n469), .IN4(n3437), .Q(n2160)
         );
  OA221X1 U1276 ( .IN1(n277), .IN2(n3434), .IN3(n309), .IN4(n3431), .IN5(n2161), .Q(n2156) );
  OA22X1 U1277 ( .IN1(n373), .IN2(n3428), .IN3(n341), .IN4(n3425), .Q(n2161)
         );
  OA222X1 U1278 ( .IN1(n181), .IN2(n3422), .IN3(n245), .IN4(n3419), .IN5(n213), 
        .IN6(n3416), .Q(n2155) );
  NAND4X0 U1279 ( .IN1(n2162), .IN2(n2163), .IN3(n2164), .IN4(n2165), .QN(
        n2153) );
  OA221X1 U1280 ( .IN1(n117), .IN2(n3413), .IN3(n85), .IN4(n3410), .IN5(n2166), 
        .Q(n2165) );
  OA22X1 U1281 ( .IN1(n149), .IN2(n3407), .IN3(n53), .IN4(n3404), .Q(n2166) );
  OA221X1 U1282 ( .IN1(n917), .IN2(n3401), .IN3(n949), .IN4(n3398), .IN5(n2167), .Q(n2164) );
  OA22X1 U1283 ( .IN1(n21), .IN2(n3395), .IN3(n981), .IN4(n3392), .Q(n2167) );
  OA221X1 U1284 ( .IN1(n789), .IN2(n3389), .IN3(n821), .IN4(n3386), .IN5(n2168), .Q(n2163) );
  OA22X1 U1285 ( .IN1(n885), .IN2(n3383), .IN3(n853), .IN4(n3380), .Q(n2168)
         );
  OA221X1 U1286 ( .IN1(n725), .IN2(n3377), .IN3(n757), .IN4(n3374), .IN5(n2169), .Q(n2162) );
  OA22X1 U1287 ( .IN1(n693), .IN2(n3371), .IN3(n661), .IN4(n3368), .Q(n2169)
         );
  OR2X1 U1288 ( .IN1(n2170), .IN2(n2171), .Q(rd_dataA[10]) );
  NAND4X0 U1289 ( .IN1(n2172), .IN2(n2173), .IN3(n2174), .IN4(n2175), .QN(
        n2171) );
  OA221X1 U1290 ( .IN1(n534), .IN2(n3458), .IN3(n566), .IN4(n3455), .IN5(n2176), .Q(n2175) );
  OA22X1 U1291 ( .IN1(n630), .IN2(n3452), .IN3(n598), .IN4(n3449), .Q(n2176)
         );
  OA221X1 U1292 ( .IN1(n406), .IN2(n3446), .IN3(n438), .IN4(n3443), .IN5(n2177), .Q(n2174) );
  OA22X1 U1293 ( .IN1(n502), .IN2(n3440), .IN3(n470), .IN4(n3437), .Q(n2177)
         );
  OA221X1 U1294 ( .IN1(n278), .IN2(n3434), .IN3(n310), .IN4(n3431), .IN5(n2178), .Q(n2173) );
  OA22X1 U1295 ( .IN1(n374), .IN2(n3428), .IN3(n342), .IN4(n3425), .Q(n2178)
         );
  OA222X1 U1296 ( .IN1(n182), .IN2(n3422), .IN3(n246), .IN4(n3419), .IN5(n214), 
        .IN6(n3416), .Q(n2172) );
  NAND4X0 U1297 ( .IN1(n2179), .IN2(n2180), .IN3(n2181), .IN4(n2182), .QN(
        n2170) );
  OA221X1 U1298 ( .IN1(n118), .IN2(n3413), .IN3(n86), .IN4(n3410), .IN5(n2183), 
        .Q(n2182) );
  OA22X1 U1299 ( .IN1(n150), .IN2(n3407), .IN3(n54), .IN4(n3404), .Q(n2183) );
  OA221X1 U1300 ( .IN1(n918), .IN2(n3401), .IN3(n950), .IN4(n3398), .IN5(n2184), .Q(n2181) );
  OA22X1 U1301 ( .IN1(n22), .IN2(n3395), .IN3(n982), .IN4(n3392), .Q(n2184) );
  OA221X1 U1302 ( .IN1(n790), .IN2(n3389), .IN3(n822), .IN4(n3386), .IN5(n2185), .Q(n2180) );
  OA22X1 U1303 ( .IN1(n886), .IN2(n3383), .IN3(n854), .IN4(n3380), .Q(n2185)
         );
  OA221X1 U1304 ( .IN1(n726), .IN2(n3377), .IN3(n758), .IN4(n3374), .IN5(n2186), .Q(n2179) );
  OA22X1 U1305 ( .IN1(n694), .IN2(n3371), .IN3(n662), .IN4(n3368), .Q(n2186)
         );
  OR2X1 U1306 ( .IN1(n2187), .IN2(n2188), .Q(rd_dataA[0]) );
  NAND4X0 U1307 ( .IN1(n2189), .IN2(n2190), .IN3(n2191), .IN4(n2192), .QN(
        n2188) );
  OA221X1 U1308 ( .IN1(n544), .IN2(n3458), .IN3(n576), .IN4(n3455), .IN5(n2193), .Q(n2192) );
  OA22X1 U1309 ( .IN1(n640), .IN2(n3452), .IN3(n608), .IN4(n3449), .Q(n2193)
         );
  OA221X1 U1310 ( .IN1(n416), .IN2(n3446), .IN3(n448), .IN4(n3443), .IN5(n2198), .Q(n2191) );
  OA22X1 U1311 ( .IN1(n512), .IN2(n3440), .IN3(n480), .IN4(n3437), .Q(n2198)
         );
  OA221X1 U1312 ( .IN1(n288), .IN2(n3434), .IN3(n320), .IN4(n3431), .IN5(n2201), .Q(n2190) );
  OA22X1 U1313 ( .IN1(n384), .IN2(n3428), .IN3(n352), .IN4(n3425), .Q(n2201)
         );
  OA222X1 U1314 ( .IN1(n192), .IN2(n3422), .IN3(n256), .IN4(n3419), .IN5(n224), 
        .IN6(n3416), .Q(n2189) );
  NAND4X0 U1315 ( .IN1(n2206), .IN2(n2207), .IN3(n2208), .IN4(n2209), .QN(
        n2187) );
  OA221X1 U1316 ( .IN1(n128), .IN2(n3413), .IN3(n96), .IN4(n3410), .IN5(n2210), 
        .Q(n2209) );
  OA22X1 U1317 ( .IN1(n160), .IN2(n3407), .IN3(n64), .IN4(n3404), .Q(n2210) );
  AND3X1 U1318 ( .IN1(rd_addrA[2]), .IN2(rd_addrA[1]), .IN3(rd_addrA[3]), .Q(
        n2195) );
  AND2X1 U1319 ( .IN1(n2213), .IN2(rd_addrA[3]), .Q(n2197) );
  OA221X1 U1320 ( .IN1(n928), .IN2(n3401), .IN3(n960), .IN4(n3398), .IN5(n2214), .Q(n2208) );
  OA22X1 U1321 ( .IN1(n32), .IN2(n3395), .IN3(n992), .IN4(n3392), .Q(n2214) );
  AND2X1 U1322 ( .IN1(n2215), .IN2(rd_addrA[1]), .Q(n2199) );
  AND2X1 U1323 ( .IN1(n2215), .IN2(n3746), .Q(n2200) );
  OA221X1 U1324 ( .IN1(n800), .IN2(n3389), .IN3(n832), .IN4(n3386), .IN5(n2216), .Q(n2207) );
  OA22X1 U1325 ( .IN1(n896), .IN2(n3383), .IN3(n864), .IN4(n3380), .Q(n2216)
         );
  AND2X1 U1326 ( .IN1(n2217), .IN2(rd_addrA[2]), .Q(n2202) );
  AND2X1 U1327 ( .IN1(n2213), .IN2(n3744), .Q(n2203) );
  OA221X1 U1328 ( .IN1(n736), .IN2(n3377), .IN3(n768), .IN4(n3374), .IN5(n2218), .Q(n2206) );
  OA22X1 U1329 ( .IN1(n704), .IN2(n3371), .IN3(n672), .IN4(n3368), .Q(n2218)
         );
  AND3X1 U1330 ( .IN1(n3745), .IN2(n3744), .IN3(n3746), .Q(n2205) );
  AND2X1 U1331 ( .IN1(n2217), .IN2(n3745), .Q(n2204) );
  AO22X1 U1332 ( .IN1(n3588), .IN2(n3363), .IN3(elem30[12]), .IN4(n2219), .Q(
        n3208) );
  AO22X1 U1333 ( .IN1(n3591), .IN2(n3365), .IN3(elem30[13]), .IN4(n3362), .Q(
        n3209) );
  AO22X1 U1334 ( .IN1(n3594), .IN2(n3365), .IN3(elem30[14]), .IN4(n2219), .Q(
        n3210) );
  AO22X1 U1335 ( .IN1(n3597), .IN2(n3365), .IN3(elem30[15]), .IN4(n2219), .Q(
        n3211) );
  AO22X1 U1336 ( .IN1(n3600), .IN2(n3365), .IN3(elem30[16]), .IN4(n2219), .Q(
        n3212) );
  AO22X1 U1337 ( .IN1(n3603), .IN2(n3364), .IN3(elem30[17]), .IN4(n2219), .Q(
        n3213) );
  AO22X1 U1338 ( .IN1(n3606), .IN2(n3363), .IN3(elem30[18]), .IN4(n2219), .Q(
        n3214) );
  AO22X1 U1339 ( .IN1(n3609), .IN2(n3365), .IN3(elem30[19]), .IN4(n2219), .Q(
        n3215) );
  AO22X1 U1340 ( .IN1(n3612), .IN2(n3364), .IN3(elem30[20]), .IN4(n3362), .Q(
        n3216) );
  AO22X1 U1341 ( .IN1(n3615), .IN2(n3363), .IN3(elem30[21]), .IN4(n3362), .Q(
        n3217) );
  AO22X1 U1342 ( .IN1(n3618), .IN2(n3365), .IN3(elem30[22]), .IN4(n3362), .Q(
        n3218) );
  AO22X1 U1343 ( .IN1(n3621), .IN2(n3363), .IN3(elem30[23]), .IN4(n3362), .Q(
        n3219) );
  AO22X1 U1344 ( .IN1(n3624), .IN2(n3363), .IN3(elem30[24]), .IN4(n3362), .Q(
        n3220) );
  AO22X1 U1345 ( .IN1(n3627), .IN2(n3363), .IN3(elem30[25]), .IN4(n3362), .Q(
        n3221) );
  AO22X1 U1346 ( .IN1(n3630), .IN2(n3363), .IN3(elem30[26]), .IN4(n3362), .Q(
        n3222) );
  AO22X1 U1347 ( .IN1(n3633), .IN2(n3363), .IN3(elem30[27]), .IN4(n3362), .Q(
        n3223) );
  AO22X1 U1348 ( .IN1(n3636), .IN2(n3363), .IN3(elem30[28]), .IN4(n3362), .Q(
        n3224) );
  AO22X1 U1349 ( .IN1(n3639), .IN2(n3363), .IN3(elem30[29]), .IN4(n3362), .Q(
        n3225) );
  AO22X1 U1350 ( .IN1(n3642), .IN2(n3364), .IN3(elem30[30]), .IN4(n3362), .Q(
        n3226) );
  AO22X1 U1351 ( .IN1(n3645), .IN2(n3364), .IN3(elem30[31]), .IN4(n3362), .Q(
        n3227) );
  AO22X1 U1352 ( .IN1(n3552), .IN2(n3360), .IN3(elem27[0]), .IN4(n3357), .Q(
        n3228) );
  AO22X1 U1353 ( .IN1(n3555), .IN2(n3360), .IN3(elem27[1]), .IN4(n2220), .Q(
        n3229) );
  AO22X1 U1354 ( .IN1(n3558), .IN2(n3360), .IN3(elem27[2]), .IN4(n2220), .Q(
        n3230) );
  AO22X1 U1355 ( .IN1(n3561), .IN2(n3360), .IN3(elem27[3]), .IN4(n2220), .Q(
        n3231) );
  AO22X1 U1356 ( .IN1(n3564), .IN2(n3360), .IN3(elem27[4]), .IN4(n2220), .Q(
        n3232) );
  AO22X1 U1357 ( .IN1(n3567), .IN2(n3360), .IN3(elem27[5]), .IN4(n2220), .Q(
        n3233) );
  AO22X1 U1358 ( .IN1(n3570), .IN2(n3360), .IN3(elem27[6]), .IN4(n2220), .Q(
        n3234) );
  AO22X1 U1359 ( .IN1(n3573), .IN2(n3359), .IN3(elem27[7]), .IN4(n2220), .Q(
        n3235) );
  AO22X1 U1360 ( .IN1(n3576), .IN2(n3359), .IN3(elem27[8]), .IN4(n3357), .Q(
        n3236) );
  AO22X1 U1361 ( .IN1(n3579), .IN2(n3359), .IN3(elem27[9]), .IN4(n3357), .Q(
        n3237) );
  AO22X1 U1362 ( .IN1(n3582), .IN2(n3359), .IN3(elem27[10]), .IN4(n3357), .Q(
        n3238) );
  AO22X1 U1363 ( .IN1(n3585), .IN2(n3359), .IN3(elem27[11]), .IN4(n3357), .Q(
        n3239) );
  AO22X1 U1364 ( .IN1(n3359), .IN2(n3588), .IN3(elem27[12]), .IN4(n3357), .Q(
        n3240) );
  AO22X1 U1365 ( .IN1(n3359), .IN2(n3591), .IN3(elem27[13]), .IN4(n3357), .Q(
        n3241) );
  AO22X1 U1366 ( .IN1(n3358), .IN2(n3594), .IN3(elem27[14]), .IN4(n3357), .Q(
        n3242) );
  AO22X1 U1367 ( .IN1(n3359), .IN2(n3597), .IN3(elem27[15]), .IN4(n3357), .Q(
        n3243) );
  AO22X1 U1368 ( .IN1(n3360), .IN2(n3600), .IN3(elem27[16]), .IN4(n3357), .Q(
        n3244) );
  AO22X1 U1369 ( .IN1(n3359), .IN2(n3603), .IN3(elem27[17]), .IN4(n3357), .Q(
        n3245) );
  AO22X1 U1370 ( .IN1(n3358), .IN2(n3606), .IN3(elem27[18]), .IN4(n3357), .Q(
        n3246) );
  AO22X1 U1371 ( .IN1(n3360), .IN2(n3609), .IN3(elem27[19]), .IN4(n3357), .Q(
        n3247) );
  AO22X1 U1372 ( .IN1(n3358), .IN2(n3612), .IN3(elem27[20]), .IN4(n3356), .Q(
        n3248) );
  AO22X1 U1373 ( .IN1(n3358), .IN2(n3615), .IN3(elem27[21]), .IN4(n3356), .Q(
        n3249) );
  AO22X1 U1374 ( .IN1(n3358), .IN2(n3618), .IN3(elem27[22]), .IN4(n3356), .Q(
        n3250) );
  AO22X1 U1375 ( .IN1(n3358), .IN2(n3621), .IN3(elem27[23]), .IN4(n3356), .Q(
        n3251) );
  AO22X1 U1376 ( .IN1(n3358), .IN2(n3624), .IN3(elem27[24]), .IN4(n3356), .Q(
        n3252) );
  AO22X1 U1377 ( .IN1(n3358), .IN2(n3627), .IN3(elem27[25]), .IN4(n3356), .Q(
        n3253) );
  AO22X1 U1378 ( .IN1(n3358), .IN2(n3630), .IN3(elem27[26]), .IN4(n3356), .Q(
        n3254) );
  AO22X1 U1379 ( .IN1(n3360), .IN2(n3633), .IN3(elem27[27]), .IN4(n3356), .Q(
        n3255) );
  AO22X1 U1380 ( .IN1(n3360), .IN2(n3636), .IN3(elem27[28]), .IN4(n3356), .Q(
        n3256) );
  AO22X1 U1381 ( .IN1(n3360), .IN2(n3639), .IN3(elem27[29]), .IN4(n3356), .Q(
        n3257) );
  AO22X1 U1382 ( .IN1(n3359), .IN2(n3642), .IN3(elem27[30]), .IN4(n3356), .Q(
        n3258) );
  AO22X1 U1383 ( .IN1(n3360), .IN2(n3645), .IN3(elem27[31]), .IN4(n3356), .Q(
        n3259) );
  AO22X1 U1384 ( .IN1(n3353), .IN2(n3552), .IN3(elem26[0]), .IN4(n2223), .Q(
        n2268) );
  AO22X1 U1385 ( .IN1(n3353), .IN2(n3555), .IN3(elem26[1]), .IN4(n2223), .Q(
        n2269) );
  AO22X1 U1386 ( .IN1(n3353), .IN2(n3558), .IN3(elem26[2]), .IN4(n2223), .Q(
        n2270) );
  AO22X1 U1387 ( .IN1(n3353), .IN2(n3561), .IN3(elem26[3]), .IN4(n2223), .Q(
        n2271) );
  AO22X1 U1388 ( .IN1(n3354), .IN2(n3564), .IN3(elem26[4]), .IN4(n2223), .Q(
        n2272) );
  AO22X1 U1389 ( .IN1(n3355), .IN2(n3567), .IN3(elem26[5]), .IN4(n2223), .Q(
        n2273) );
  AO22X1 U1390 ( .IN1(n3355), .IN2(n3570), .IN3(elem26[6]), .IN4(n2223), .Q(
        n2274) );
  AO22X1 U1391 ( .IN1(n3354), .IN2(n3573), .IN3(elem26[7]), .IN4(n2223), .Q(
        n2275) );
  AO22X1 U1392 ( .IN1(n3355), .IN2(n3576), .IN3(elem26[8]), .IN4(n3352), .Q(
        n2276) );
  AO22X1 U1393 ( .IN1(n3355), .IN2(n3579), .IN3(elem26[9]), .IN4(n3352), .Q(
        n2277) );
  AO22X1 U1394 ( .IN1(n3354), .IN2(n3582), .IN3(elem26[10]), .IN4(n3352), .Q(
        n2278) );
  AO22X1 U1395 ( .IN1(n3354), .IN2(n3585), .IN3(elem26[11]), .IN4(n3352), .Q(
        n2279) );
  AO22X1 U1396 ( .IN1(n3354), .IN2(n3588), .IN3(elem26[12]), .IN4(n3352), .Q(
        n2280) );
  AO22X1 U1397 ( .IN1(n3354), .IN2(n3591), .IN3(elem26[13]), .IN4(n3352), .Q(
        n2281) );
  AO22X1 U1398 ( .IN1(n3354), .IN2(n3594), .IN3(elem26[14]), .IN4(n3352), .Q(
        n2282) );
  AO22X1 U1399 ( .IN1(n3354), .IN2(n3597), .IN3(elem26[15]), .IN4(n3352), .Q(
        n2283) );
  AO22X1 U1400 ( .IN1(n3354), .IN2(n3600), .IN3(elem26[16]), .IN4(n3352), .Q(
        n2284) );
  AO22X1 U1401 ( .IN1(n3354), .IN2(n3603), .IN3(elem26[17]), .IN4(n3352), .Q(
        n2285) );
  AO22X1 U1402 ( .IN1(n3354), .IN2(n3606), .IN3(elem26[18]), .IN4(n3352), .Q(
        n2286) );
  AO22X1 U1403 ( .IN1(n3355), .IN2(n3609), .IN3(elem26[19]), .IN4(n3352), .Q(
        n2287) );
  AO22X1 U1404 ( .IN1(n3354), .IN2(n3612), .IN3(elem26[20]), .IN4(n3351), .Q(
        n2288) );
  AO22X1 U1405 ( .IN1(n3355), .IN2(n3615), .IN3(elem26[21]), .IN4(n3351), .Q(
        n2289) );
  AO22X1 U1406 ( .IN1(n3354), .IN2(n3618), .IN3(elem26[22]), .IN4(n3351), .Q(
        n2290) );
  AO22X1 U1407 ( .IN1(n3355), .IN2(n3621), .IN3(elem26[23]), .IN4(n3351), .Q(
        n2291) );
  AO22X1 U1408 ( .IN1(n3354), .IN2(n3624), .IN3(elem26[24]), .IN4(n3351), .Q(
        n2292) );
  AO22X1 U1409 ( .IN1(n3355), .IN2(n3627), .IN3(elem26[25]), .IN4(n3351), .Q(
        n2293) );
  AO22X1 U1410 ( .IN1(n3355), .IN2(n3630), .IN3(elem26[26]), .IN4(n3351), .Q(
        n2294) );
  AO22X1 U1411 ( .IN1(n3355), .IN2(n3633), .IN3(elem26[27]), .IN4(n3351), .Q(
        n2295) );
  AO22X1 U1412 ( .IN1(n3355), .IN2(n3636), .IN3(elem26[28]), .IN4(n3351), .Q(
        n2296) );
  AO22X1 U1413 ( .IN1(n3355), .IN2(n3639), .IN3(elem26[29]), .IN4(n3351), .Q(
        n2297) );
  AO22X1 U1414 ( .IN1(n3355), .IN2(n3642), .IN3(elem26[30]), .IN4(n3351), .Q(
        n2298) );
  AO22X1 U1415 ( .IN1(n3355), .IN2(n3645), .IN3(elem26[31]), .IN4(n3351), .Q(
        n2299) );
  AO22X1 U1416 ( .IN1(n3349), .IN2(n3554), .IN3(elem25[0]), .IN4(n2225), .Q(
        n2300) );
  AO22X1 U1417 ( .IN1(n3348), .IN2(n3557), .IN3(elem25[1]), .IN4(n3347), .Q(
        n2301) );
  AO22X1 U1418 ( .IN1(n3348), .IN2(n3560), .IN3(elem25[2]), .IN4(n2225), .Q(
        n2302) );
  AO22X1 U1419 ( .IN1(n3348), .IN2(n3563), .IN3(elem25[3]), .IN4(n2225), .Q(
        n2303) );
  AO22X1 U1420 ( .IN1(n3348), .IN2(n3566), .IN3(elem25[4]), .IN4(n2225), .Q(
        n2304) );
  AO22X1 U1421 ( .IN1(n3350), .IN2(n3569), .IN3(elem25[5]), .IN4(n2225), .Q(
        n2305) );
  AO22X1 U1422 ( .IN1(n3349), .IN2(n3572), .IN3(elem25[6]), .IN4(n2225), .Q(
        n2306) );
  AO22X1 U1423 ( .IN1(n3348), .IN2(n3575), .IN3(elem25[7]), .IN4(n2225), .Q(
        n2307) );
  AO22X1 U1424 ( .IN1(n3350), .IN2(n3578), .IN3(elem25[8]), .IN4(n3347), .Q(
        n2308) );
  AO22X1 U1425 ( .IN1(n3349), .IN2(n3581), .IN3(elem25[9]), .IN4(n3347), .Q(
        n2309) );
  AO22X1 U1426 ( .IN1(n3348), .IN2(n3584), .IN3(elem25[10]), .IN4(n3347), .Q(
        n2310) );
  AO22X1 U1427 ( .IN1(n3348), .IN2(n3587), .IN3(elem25[11]), .IN4(n3347), .Q(
        n2311) );
  AO22X1 U1428 ( .IN1(n3348), .IN2(n3588), .IN3(elem25[12]), .IN4(n3347), .Q(
        n2312) );
  AO22X1 U1429 ( .IN1(n3348), .IN2(n3591), .IN3(elem25[13]), .IN4(n3347), .Q(
        n2313) );
  AO22X1 U1430 ( .IN1(n3348), .IN2(n3594), .IN3(elem25[14]), .IN4(n3347), .Q(
        n2314) );
  AO22X1 U1431 ( .IN1(n3348), .IN2(n3597), .IN3(elem25[15]), .IN4(n3347), .Q(
        n2315) );
  AO22X1 U1432 ( .IN1(n3348), .IN2(n3600), .IN3(elem25[16]), .IN4(n3347), .Q(
        n2316) );
  AO22X1 U1433 ( .IN1(n3348), .IN2(n3603), .IN3(elem25[17]), .IN4(n3347), .Q(
        n2317) );
  AO22X1 U1434 ( .IN1(n3349), .IN2(n3606), .IN3(elem25[18]), .IN4(n3347), .Q(
        n2318) );
  AO22X1 U1435 ( .IN1(n3349), .IN2(n3609), .IN3(elem25[19]), .IN4(n3347), .Q(
        n2319) );
  AO22X1 U1436 ( .IN1(n3349), .IN2(n3612), .IN3(elem25[20]), .IN4(n3346), .Q(
        n2320) );
  AO22X1 U1437 ( .IN1(n3349), .IN2(n3615), .IN3(elem25[21]), .IN4(n3346), .Q(
        n2321) );
  AO22X1 U1438 ( .IN1(n3349), .IN2(n3618), .IN3(elem25[22]), .IN4(n3346), .Q(
        n2322) );
  AO22X1 U1439 ( .IN1(n3349), .IN2(n3621), .IN3(elem25[23]), .IN4(n3346), .Q(
        n2323) );
  AO22X1 U1440 ( .IN1(n3349), .IN2(n3624), .IN3(elem25[24]), .IN4(n3346), .Q(
        n2324) );
  AO22X1 U1441 ( .IN1(n3350), .IN2(n3627), .IN3(elem25[25]), .IN4(n3346), .Q(
        n2325) );
  AO22X1 U1442 ( .IN1(n3350), .IN2(n3630), .IN3(elem25[26]), .IN4(n3346), .Q(
        n2326) );
  AO22X1 U1443 ( .IN1(n3350), .IN2(n3633), .IN3(elem25[27]), .IN4(n3346), .Q(
        n2327) );
  AO22X1 U1444 ( .IN1(n3350), .IN2(n3636), .IN3(elem25[28]), .IN4(n3346), .Q(
        n2328) );
  AO22X1 U1445 ( .IN1(n3350), .IN2(n3639), .IN3(elem25[29]), .IN4(n3346), .Q(
        n2329) );
  AO22X1 U1446 ( .IN1(n3350), .IN2(n3642), .IN3(elem25[30]), .IN4(n3346), .Q(
        n2330) );
  AO22X1 U1447 ( .IN1(n3350), .IN2(n3645), .IN3(elem25[31]), .IN4(n3346), .Q(
        n2331) );
  AO22X1 U1448 ( .IN1(n3344), .IN2(n3554), .IN3(elem24[0]), .IN4(n2227), .Q(
        n2332) );
  AO22X1 U1449 ( .IN1(n3343), .IN2(n3557), .IN3(elem24[1]), .IN4(n3342), .Q(
        n2333) );
  AO22X1 U1450 ( .IN1(n3343), .IN2(n3560), .IN3(elem24[2]), .IN4(n2227), .Q(
        n2334) );
  AO22X1 U1451 ( .IN1(n3343), .IN2(n3563), .IN3(elem24[3]), .IN4(n2227), .Q(
        n2335) );
  AO22X1 U1452 ( .IN1(n3343), .IN2(n3566), .IN3(elem24[4]), .IN4(n2227), .Q(
        n2336) );
  AO22X1 U1453 ( .IN1(n3345), .IN2(n3569), .IN3(elem24[5]), .IN4(n2227), .Q(
        n2337) );
  AO22X1 U1454 ( .IN1(n3344), .IN2(n3572), .IN3(elem24[6]), .IN4(n2227), .Q(
        n2338) );
  AO22X1 U1455 ( .IN1(n3343), .IN2(n3575), .IN3(elem24[7]), .IN4(n2227), .Q(
        n2339) );
  AO22X1 U1456 ( .IN1(n3345), .IN2(n3578), .IN3(elem24[8]), .IN4(n3342), .Q(
        n2340) );
  AO22X1 U1457 ( .IN1(n3344), .IN2(n3581), .IN3(elem24[9]), .IN4(n3342), .Q(
        n2341) );
  AO22X1 U1458 ( .IN1(n3343), .IN2(n3584), .IN3(elem24[10]), .IN4(n3342), .Q(
        n2342) );
  AO22X1 U1459 ( .IN1(n3343), .IN2(n3587), .IN3(elem24[11]), .IN4(n3342), .Q(
        n2343) );
  AO22X1 U1460 ( .IN1(n3343), .IN2(n3588), .IN3(elem24[12]), .IN4(n3342), .Q(
        n2344) );
  AO22X1 U1461 ( .IN1(n3343), .IN2(n3591), .IN3(elem24[13]), .IN4(n3342), .Q(
        n2345) );
  AO22X1 U1462 ( .IN1(n3343), .IN2(n3594), .IN3(elem24[14]), .IN4(n3342), .Q(
        n2346) );
  AO22X1 U1463 ( .IN1(n3343), .IN2(n3597), .IN3(elem24[15]), .IN4(n3342), .Q(
        n2347) );
  AO22X1 U1464 ( .IN1(n3343), .IN2(n3600), .IN3(elem24[16]), .IN4(n3342), .Q(
        n2348) );
  AO22X1 U1465 ( .IN1(n3343), .IN2(n3603), .IN3(elem24[17]), .IN4(n3342), .Q(
        n2349) );
  AO22X1 U1466 ( .IN1(n3344), .IN2(n3606), .IN3(elem24[18]), .IN4(n3342), .Q(
        n2350) );
  AO22X1 U1467 ( .IN1(n3344), .IN2(n3609), .IN3(elem24[19]), .IN4(n3342), .Q(
        n2351) );
  AO22X1 U1468 ( .IN1(n3344), .IN2(n3612), .IN3(elem24[20]), .IN4(n3341), .Q(
        n2352) );
  AO22X1 U1469 ( .IN1(n3344), .IN2(n3615), .IN3(elem24[21]), .IN4(n3341), .Q(
        n2353) );
  AO22X1 U1470 ( .IN1(n3344), .IN2(n3618), .IN3(elem24[22]), .IN4(n3341), .Q(
        n2354) );
  AO22X1 U1471 ( .IN1(n3344), .IN2(n3621), .IN3(elem24[23]), .IN4(n3341), .Q(
        n2355) );
  AO22X1 U1472 ( .IN1(n3344), .IN2(n3624), .IN3(elem24[24]), .IN4(n3341), .Q(
        n2356) );
  AO22X1 U1473 ( .IN1(n3345), .IN2(n3627), .IN3(elem24[25]), .IN4(n3341), .Q(
        n2357) );
  AO22X1 U1474 ( .IN1(n3345), .IN2(n3630), .IN3(elem24[26]), .IN4(n3341), .Q(
        n2358) );
  AO22X1 U1475 ( .IN1(n3345), .IN2(n3633), .IN3(elem24[27]), .IN4(n3341), .Q(
        n2359) );
  AO22X1 U1476 ( .IN1(n3345), .IN2(n3636), .IN3(elem24[28]), .IN4(n3341), .Q(
        n2360) );
  AO22X1 U1477 ( .IN1(n3345), .IN2(n3639), .IN3(elem24[29]), .IN4(n3341), .Q(
        n2361) );
  AO22X1 U1478 ( .IN1(n3345), .IN2(n3642), .IN3(elem24[30]), .IN4(n3341), .Q(
        n2362) );
  AO22X1 U1479 ( .IN1(n3345), .IN2(n3645), .IN3(elem24[31]), .IN4(n3341), .Q(
        n2363) );
  AND2X1 U1480 ( .IN1(n2229), .IN2(n2230), .Q(n2222) );
  AO22X1 U1481 ( .IN1(n3338), .IN2(n3554), .IN3(elem23[0]), .IN4(n2231), .Q(
        n2364) );
  AO22X1 U1482 ( .IN1(n3338), .IN2(n3557), .IN3(elem23[1]), .IN4(n2231), .Q(
        n2365) );
  AO22X1 U1483 ( .IN1(n3338), .IN2(n3560), .IN3(elem23[2]), .IN4(n2231), .Q(
        n2366) );
  AO22X1 U1484 ( .IN1(n3338), .IN2(n3563), .IN3(elem23[3]), .IN4(n2231), .Q(
        n2367) );
  AO22X1 U1485 ( .IN1(n3339), .IN2(n3566), .IN3(elem23[4]), .IN4(n2231), .Q(
        n2368) );
  AO22X1 U1486 ( .IN1(n3340), .IN2(n3569), .IN3(elem23[5]), .IN4(n2231), .Q(
        n2369) );
  AO22X1 U1487 ( .IN1(n3340), .IN2(n3572), .IN3(elem23[6]), .IN4(n2231), .Q(
        n2370) );
  AO22X1 U1488 ( .IN1(n3339), .IN2(n3575), .IN3(elem23[7]), .IN4(n2231), .Q(
        n2371) );
  AO22X1 U1489 ( .IN1(n3340), .IN2(n3578), .IN3(elem23[8]), .IN4(n3337), .Q(
        n2372) );
  AO22X1 U1490 ( .IN1(n3340), .IN2(n3581), .IN3(elem23[9]), .IN4(n3337), .Q(
        n2373) );
  AO22X1 U1491 ( .IN1(n3339), .IN2(n3584), .IN3(elem23[10]), .IN4(n3337), .Q(
        n2374) );
  AO22X1 U1492 ( .IN1(n3339), .IN2(n3587), .IN3(elem23[11]), .IN4(n3337), .Q(
        n2375) );
  AO22X1 U1493 ( .IN1(n3339), .IN2(n3588), .IN3(elem23[12]), .IN4(n3337), .Q(
        n2376) );
  AO22X1 U1494 ( .IN1(n3339), .IN2(n3591), .IN3(elem23[13]), .IN4(n3337), .Q(
        n2377) );
  AO22X1 U1495 ( .IN1(n3339), .IN2(n3594), .IN3(elem23[14]), .IN4(n3337), .Q(
        n2378) );
  AO22X1 U1496 ( .IN1(n3339), .IN2(n3597), .IN3(elem23[15]), .IN4(n3337), .Q(
        n2379) );
  AO22X1 U1497 ( .IN1(n3339), .IN2(n3600), .IN3(elem23[16]), .IN4(n3337), .Q(
        n2380) );
  AO22X1 U1498 ( .IN1(n3339), .IN2(n3603), .IN3(elem23[17]), .IN4(n3337), .Q(
        n2381) );
  AO22X1 U1499 ( .IN1(n3339), .IN2(n3606), .IN3(elem23[18]), .IN4(n3337), .Q(
        n2382) );
  AO22X1 U1500 ( .IN1(n3340), .IN2(n3609), .IN3(elem23[19]), .IN4(n3337), .Q(
        n2383) );
  AO22X1 U1501 ( .IN1(n3339), .IN2(n3612), .IN3(elem23[20]), .IN4(n3336), .Q(
        n2384) );
  AO22X1 U1502 ( .IN1(n3340), .IN2(n3615), .IN3(elem23[21]), .IN4(n3336), .Q(
        n2385) );
  AO22X1 U1503 ( .IN1(n3339), .IN2(n3618), .IN3(elem23[22]), .IN4(n3336), .Q(
        n2386) );
  AO22X1 U1504 ( .IN1(n3340), .IN2(n3621), .IN3(elem23[23]), .IN4(n3336), .Q(
        n2387) );
  AO22X1 U1505 ( .IN1(n3339), .IN2(n3624), .IN3(elem23[24]), .IN4(n3336), .Q(
        n2388) );
  AO22X1 U1506 ( .IN1(n3340), .IN2(n3627), .IN3(elem23[25]), .IN4(n3336), .Q(
        n2389) );
  AO22X1 U1507 ( .IN1(n3340), .IN2(n3630), .IN3(elem23[26]), .IN4(n3336), .Q(
        n2390) );
  AO22X1 U1508 ( .IN1(n3340), .IN2(n3633), .IN3(elem23[27]), .IN4(n3336), .Q(
        n2391) );
  AO22X1 U1509 ( .IN1(n3340), .IN2(n3636), .IN3(elem23[28]), .IN4(n3336), .Q(
        n2392) );
  AO22X1 U1510 ( .IN1(n3340), .IN2(n3639), .IN3(elem23[29]), .IN4(n3336), .Q(
        n2393) );
  AO22X1 U1511 ( .IN1(n3340), .IN2(n3642), .IN3(elem23[30]), .IN4(n3336), .Q(
        n2394) );
  AO22X1 U1512 ( .IN1(n3340), .IN2(n3645), .IN3(elem23[31]), .IN4(n3336), .Q(
        n2395) );
  AO22X1 U1513 ( .IN1(n3333), .IN2(n3554), .IN3(elem22[0]), .IN4(n2233), .Q(
        n2396) );
  AO22X1 U1514 ( .IN1(n3333), .IN2(n3557), .IN3(elem22[1]), .IN4(n2233), .Q(
        n2397) );
  AO22X1 U1515 ( .IN1(n3333), .IN2(n3560), .IN3(elem22[2]), .IN4(n2233), .Q(
        n2398) );
  AO22X1 U1516 ( .IN1(n3333), .IN2(n3563), .IN3(elem22[3]), .IN4(n2233), .Q(
        n2399) );
  AO22X1 U1517 ( .IN1(n3334), .IN2(n3566), .IN3(elem22[4]), .IN4(n2233), .Q(
        n2400) );
  AO22X1 U1518 ( .IN1(n3335), .IN2(n3569), .IN3(elem22[5]), .IN4(n2233), .Q(
        n2401) );
  AO22X1 U1519 ( .IN1(n3335), .IN2(n3572), .IN3(elem22[6]), .IN4(n2233), .Q(
        n2402) );
  AO22X1 U1520 ( .IN1(n3334), .IN2(n3575), .IN3(elem22[7]), .IN4(n2233), .Q(
        n2403) );
  AO22X1 U1521 ( .IN1(n3335), .IN2(n3578), .IN3(elem22[8]), .IN4(n3332), .Q(
        n2404) );
  AO22X1 U1522 ( .IN1(n3335), .IN2(n3581), .IN3(elem22[9]), .IN4(n3332), .Q(
        n2405) );
  AO22X1 U1523 ( .IN1(n3334), .IN2(n3584), .IN3(elem22[10]), .IN4(n3332), .Q(
        n2406) );
  AO22X1 U1524 ( .IN1(n3334), .IN2(n3587), .IN3(elem22[11]), .IN4(n3332), .Q(
        n2407) );
  AO22X1 U1525 ( .IN1(n3334), .IN2(n3588), .IN3(elem22[12]), .IN4(n3332), .Q(
        n2408) );
  AO22X1 U1526 ( .IN1(n3334), .IN2(n3591), .IN3(elem22[13]), .IN4(n3332), .Q(
        n2409) );
  AO22X1 U1527 ( .IN1(n3334), .IN2(n3594), .IN3(elem22[14]), .IN4(n3332), .Q(
        n2410) );
  AO22X1 U1528 ( .IN1(n3334), .IN2(n3597), .IN3(elem22[15]), .IN4(n3332), .Q(
        n2411) );
  AO22X1 U1529 ( .IN1(n3334), .IN2(n3600), .IN3(elem22[16]), .IN4(n3332), .Q(
        n2412) );
  AO22X1 U1530 ( .IN1(n3334), .IN2(n3603), .IN3(elem22[17]), .IN4(n3332), .Q(
        n2413) );
  AO22X1 U1531 ( .IN1(n3334), .IN2(n3606), .IN3(elem22[18]), .IN4(n3332), .Q(
        n2414) );
  AO22X1 U1532 ( .IN1(n3335), .IN2(n3609), .IN3(elem22[19]), .IN4(n3332), .Q(
        n2415) );
  AO22X1 U1533 ( .IN1(n3334), .IN2(n3612), .IN3(elem22[20]), .IN4(n3331), .Q(
        n2416) );
  AO22X1 U1534 ( .IN1(n3335), .IN2(n3615), .IN3(elem22[21]), .IN4(n3331), .Q(
        n2417) );
  AO22X1 U1535 ( .IN1(n3334), .IN2(n3618), .IN3(elem22[22]), .IN4(n3331), .Q(
        n2418) );
  AO22X1 U1536 ( .IN1(n3335), .IN2(n3621), .IN3(elem22[23]), .IN4(n3331), .Q(
        n2419) );
  AO22X1 U1537 ( .IN1(n3334), .IN2(n3624), .IN3(elem22[24]), .IN4(n3331), .Q(
        n2420) );
  AO22X1 U1538 ( .IN1(n3335), .IN2(n3627), .IN3(elem22[25]), .IN4(n3331), .Q(
        n2421) );
  AO22X1 U1539 ( .IN1(n3335), .IN2(n3630), .IN3(elem22[26]), .IN4(n3331), .Q(
        n2422) );
  AO22X1 U1540 ( .IN1(n3335), .IN2(n3633), .IN3(elem22[27]), .IN4(n3331), .Q(
        n2423) );
  AO22X1 U1541 ( .IN1(n3335), .IN2(n3636), .IN3(elem22[28]), .IN4(n3331), .Q(
        n2424) );
  AO22X1 U1542 ( .IN1(n3335), .IN2(n3639), .IN3(elem22[29]), .IN4(n3331), .Q(
        n2425) );
  AO22X1 U1543 ( .IN1(n3335), .IN2(n3642), .IN3(elem22[30]), .IN4(n3331), .Q(
        n2426) );
  AO22X1 U1544 ( .IN1(n3335), .IN2(n3645), .IN3(elem22[31]), .IN4(n3331), .Q(
        n2427) );
  AO22X1 U1545 ( .IN1(n3328), .IN2(n3554), .IN3(elem21[0]), .IN4(n2234), .Q(
        n2428) );
  AO22X1 U1546 ( .IN1(n3328), .IN2(n3557), .IN3(elem21[1]), .IN4(n2234), .Q(
        n2429) );
  AO22X1 U1547 ( .IN1(n3328), .IN2(n3560), .IN3(elem21[2]), .IN4(n2234), .Q(
        n2430) );
  AO22X1 U1548 ( .IN1(n3328), .IN2(n3563), .IN3(elem21[3]), .IN4(n2234), .Q(
        n2431) );
  AO22X1 U1549 ( .IN1(n3329), .IN2(n3566), .IN3(elem21[4]), .IN4(n2234), .Q(
        n2432) );
  AO22X1 U1550 ( .IN1(n3330), .IN2(n3569), .IN3(elem21[5]), .IN4(n2234), .Q(
        n2433) );
  AO22X1 U1551 ( .IN1(n3330), .IN2(n3572), .IN3(elem21[6]), .IN4(n2234), .Q(
        n2434) );
  AO22X1 U1552 ( .IN1(n3329), .IN2(n3575), .IN3(elem21[7]), .IN4(n2234), .Q(
        n2435) );
  AO22X1 U1553 ( .IN1(n3330), .IN2(n3578), .IN3(elem21[8]), .IN4(n3327), .Q(
        n2436) );
  AO22X1 U1554 ( .IN1(n3330), .IN2(n3581), .IN3(elem21[9]), .IN4(n3327), .Q(
        n2437) );
  AO22X1 U1555 ( .IN1(n3329), .IN2(n3584), .IN3(elem21[10]), .IN4(n3327), .Q(
        n2438) );
  AO22X1 U1556 ( .IN1(n3329), .IN2(n3587), .IN3(elem21[11]), .IN4(n3327), .Q(
        n2439) );
  AO22X1 U1557 ( .IN1(n3329), .IN2(n3588), .IN3(elem21[12]), .IN4(n3327), .Q(
        n2440) );
  AO22X1 U1558 ( .IN1(n3329), .IN2(n3591), .IN3(elem21[13]), .IN4(n3327), .Q(
        n2441) );
  AO22X1 U1559 ( .IN1(n3329), .IN2(n3594), .IN3(elem21[14]), .IN4(n3327), .Q(
        n2442) );
  AO22X1 U1560 ( .IN1(n3329), .IN2(n3597), .IN3(elem21[15]), .IN4(n3327), .Q(
        n2443) );
  AO22X1 U1561 ( .IN1(n3329), .IN2(n3600), .IN3(elem21[16]), .IN4(n3327), .Q(
        n2444) );
  AO22X1 U1562 ( .IN1(n3329), .IN2(n3603), .IN3(elem21[17]), .IN4(n3327), .Q(
        n2445) );
  AO22X1 U1563 ( .IN1(n3329), .IN2(n3606), .IN3(elem21[18]), .IN4(n3327), .Q(
        n2446) );
  AO22X1 U1564 ( .IN1(n3330), .IN2(n3609), .IN3(elem21[19]), .IN4(n3327), .Q(
        n2447) );
  AO22X1 U1565 ( .IN1(n3329), .IN2(n3612), .IN3(elem21[20]), .IN4(n3326), .Q(
        n2448) );
  AO22X1 U1566 ( .IN1(n3330), .IN2(n3615), .IN3(elem21[21]), .IN4(n3326), .Q(
        n2449) );
  AO22X1 U1567 ( .IN1(n3329), .IN2(n3618), .IN3(elem21[22]), .IN4(n3326), .Q(
        n2450) );
  AO22X1 U1568 ( .IN1(n3330), .IN2(n3621), .IN3(elem21[23]), .IN4(n3326), .Q(
        n2451) );
  AO22X1 U1569 ( .IN1(n3329), .IN2(n3624), .IN3(elem21[24]), .IN4(n3326), .Q(
        n2452) );
  AO22X1 U1570 ( .IN1(n3330), .IN2(n3627), .IN3(elem21[25]), .IN4(n3326), .Q(
        n2453) );
  AO22X1 U1571 ( .IN1(n3330), .IN2(n3630), .IN3(elem21[26]), .IN4(n3326), .Q(
        n2454) );
  AO22X1 U1572 ( .IN1(n3330), .IN2(n3633), .IN3(elem21[27]), .IN4(n3326), .Q(
        n2455) );
  AO22X1 U1573 ( .IN1(n3330), .IN2(n3636), .IN3(elem21[28]), .IN4(n3326), .Q(
        n2456) );
  AO22X1 U1574 ( .IN1(n3330), .IN2(n3639), .IN3(elem21[29]), .IN4(n3326), .Q(
        n2457) );
  AO22X1 U1575 ( .IN1(n3330), .IN2(n3642), .IN3(elem21[30]), .IN4(n3326), .Q(
        n2458) );
  AO22X1 U1576 ( .IN1(n3330), .IN2(n3645), .IN3(elem21[31]), .IN4(n3326), .Q(
        n2459) );
  AO22X1 U1577 ( .IN1(n3323), .IN2(n3554), .IN3(elem20[0]), .IN4(n2235), .Q(
        n2460) );
  AO22X1 U1578 ( .IN1(n3323), .IN2(n3557), .IN3(elem20[1]), .IN4(n2235), .Q(
        n2461) );
  AO22X1 U1579 ( .IN1(n3323), .IN2(n3560), .IN3(elem20[2]), .IN4(n2235), .Q(
        n2462) );
  AO22X1 U1580 ( .IN1(n3323), .IN2(n3563), .IN3(elem20[3]), .IN4(n2235), .Q(
        n2463) );
  AO22X1 U1581 ( .IN1(n3324), .IN2(n3566), .IN3(elem20[4]), .IN4(n2235), .Q(
        n2464) );
  AO22X1 U1582 ( .IN1(n3325), .IN2(n3569), .IN3(elem20[5]), .IN4(n2235), .Q(
        n2465) );
  AO22X1 U1583 ( .IN1(n3325), .IN2(n3572), .IN3(elem20[6]), .IN4(n2235), .Q(
        n2466) );
  AO22X1 U1584 ( .IN1(n3324), .IN2(n3575), .IN3(elem20[7]), .IN4(n2235), .Q(
        n2467) );
  AO22X1 U1585 ( .IN1(n3325), .IN2(n3578), .IN3(elem20[8]), .IN4(n3322), .Q(
        n2468) );
  AO22X1 U1586 ( .IN1(n3325), .IN2(n3581), .IN3(elem20[9]), .IN4(n3322), .Q(
        n2469) );
  AO22X1 U1587 ( .IN1(n3324), .IN2(n3584), .IN3(elem20[10]), .IN4(n3322), .Q(
        n2470) );
  AO22X1 U1588 ( .IN1(n3324), .IN2(n3587), .IN3(elem20[11]), .IN4(n3322), .Q(
        n2471) );
  AO22X1 U1589 ( .IN1(n3324), .IN2(n3588), .IN3(elem20[12]), .IN4(n3322), .Q(
        n2472) );
  AO22X1 U1590 ( .IN1(n3324), .IN2(n3591), .IN3(elem20[13]), .IN4(n3322), .Q(
        n2473) );
  AO22X1 U1591 ( .IN1(n3324), .IN2(n3594), .IN3(elem20[14]), .IN4(n3322), .Q(
        n2474) );
  AO22X1 U1592 ( .IN1(n3324), .IN2(n3597), .IN3(elem20[15]), .IN4(n3322), .Q(
        n2475) );
  AO22X1 U1593 ( .IN1(n3324), .IN2(n3600), .IN3(elem20[16]), .IN4(n3322), .Q(
        n2476) );
  AO22X1 U1594 ( .IN1(n3324), .IN2(n3603), .IN3(elem20[17]), .IN4(n3322), .Q(
        n2477) );
  AO22X1 U1595 ( .IN1(n3324), .IN2(n3606), .IN3(elem20[18]), .IN4(n3322), .Q(
        n2478) );
  AO22X1 U1596 ( .IN1(n3325), .IN2(n3609), .IN3(elem20[19]), .IN4(n3322), .Q(
        n2479) );
  AO22X1 U1597 ( .IN1(n3324), .IN2(n3612), .IN3(elem20[20]), .IN4(n3321), .Q(
        n2480) );
  AO22X1 U1598 ( .IN1(n3325), .IN2(n3615), .IN3(elem20[21]), .IN4(n3321), .Q(
        n2481) );
  AO22X1 U1599 ( .IN1(n3324), .IN2(n3618), .IN3(elem20[22]), .IN4(n3321), .Q(
        n2482) );
  AO22X1 U1600 ( .IN1(n3325), .IN2(n3621), .IN3(elem20[23]), .IN4(n3321), .Q(
        n2483) );
  AO22X1 U1601 ( .IN1(n3324), .IN2(n3624), .IN3(elem20[24]), .IN4(n3321), .Q(
        n2484) );
  AO22X1 U1602 ( .IN1(n3325), .IN2(n3627), .IN3(elem20[25]), .IN4(n3321), .Q(
        n2485) );
  AO22X1 U1603 ( .IN1(n3325), .IN2(n3630), .IN3(elem20[26]), .IN4(n3321), .Q(
        n2486) );
  AO22X1 U1604 ( .IN1(n3325), .IN2(n3633), .IN3(elem20[27]), .IN4(n3321), .Q(
        n2487) );
  AO22X1 U1605 ( .IN1(n3325), .IN2(n3636), .IN3(elem20[28]), .IN4(n3321), .Q(
        n2488) );
  AO22X1 U1606 ( .IN1(n3325), .IN2(n3639), .IN3(elem20[29]), .IN4(n3321), .Q(
        n2489) );
  AO22X1 U1607 ( .IN1(n3325), .IN2(n3642), .IN3(elem20[30]), .IN4(n3321), .Q(
        n2490) );
  AO22X1 U1608 ( .IN1(n3325), .IN2(n3645), .IN3(elem20[31]), .IN4(n3321), .Q(
        n2491) );
  AND2X1 U1609 ( .IN1(n2236), .IN2(n2230), .Q(n2232) );
  AO22X1 U1610 ( .IN1(n3318), .IN2(n3554), .IN3(elem19[0]), .IN4(n2237), .Q(
        n2492) );
  AO22X1 U1611 ( .IN1(n3318), .IN2(n3557), .IN3(elem19[1]), .IN4(n2237), .Q(
        n2493) );
  AO22X1 U1612 ( .IN1(n3318), .IN2(n3560), .IN3(elem19[2]), .IN4(n2237), .Q(
        n2494) );
  AO22X1 U1613 ( .IN1(n3318), .IN2(n3563), .IN3(elem19[3]), .IN4(n2237), .Q(
        n2495) );
  AO22X1 U1614 ( .IN1(n3319), .IN2(n3566), .IN3(elem19[4]), .IN4(n2237), .Q(
        n2496) );
  AO22X1 U1615 ( .IN1(n3320), .IN2(n3569), .IN3(elem19[5]), .IN4(n2237), .Q(
        n2497) );
  AO22X1 U1616 ( .IN1(n3320), .IN2(n3572), .IN3(elem19[6]), .IN4(n2237), .Q(
        n2498) );
  AO22X1 U1617 ( .IN1(n3319), .IN2(n3575), .IN3(elem19[7]), .IN4(n2237), .Q(
        n2499) );
  AO22X1 U1618 ( .IN1(n3320), .IN2(n3578), .IN3(elem19[8]), .IN4(n3317), .Q(
        n2500) );
  AO22X1 U1619 ( .IN1(n3320), .IN2(n3581), .IN3(elem19[9]), .IN4(n3317), .Q(
        n2501) );
  AO22X1 U1620 ( .IN1(n3319), .IN2(n3584), .IN3(elem19[10]), .IN4(n3317), .Q(
        n2502) );
  AO22X1 U1621 ( .IN1(n3319), .IN2(n3587), .IN3(elem19[11]), .IN4(n3317), .Q(
        n2503) );
  AO22X1 U1622 ( .IN1(n3319), .IN2(n3588), .IN3(elem19[12]), .IN4(n3317), .Q(
        n2504) );
  AO22X1 U1623 ( .IN1(n3319), .IN2(n3591), .IN3(elem19[13]), .IN4(n3317), .Q(
        n2505) );
  AO22X1 U1624 ( .IN1(n3319), .IN2(n3594), .IN3(elem19[14]), .IN4(n3317), .Q(
        n2506) );
  AO22X1 U1625 ( .IN1(n3319), .IN2(n3597), .IN3(elem19[15]), .IN4(n3317), .Q(
        n2507) );
  AO22X1 U1626 ( .IN1(n3319), .IN2(n3600), .IN3(elem19[16]), .IN4(n3317), .Q(
        n2508) );
  AO22X1 U1627 ( .IN1(n3319), .IN2(n3603), .IN3(elem19[17]), .IN4(n3317), .Q(
        n2509) );
  AO22X1 U1628 ( .IN1(n3319), .IN2(n3606), .IN3(elem19[18]), .IN4(n3317), .Q(
        n2510) );
  AO22X1 U1629 ( .IN1(n3320), .IN2(n3609), .IN3(elem19[19]), .IN4(n3317), .Q(
        n2511) );
  AO22X1 U1630 ( .IN1(n3319), .IN2(n3612), .IN3(elem19[20]), .IN4(n3316), .Q(
        n2512) );
  AO22X1 U1631 ( .IN1(n3320), .IN2(n3615), .IN3(elem19[21]), .IN4(n3316), .Q(
        n2513) );
  AO22X1 U1632 ( .IN1(n3319), .IN2(n3618), .IN3(elem19[22]), .IN4(n3316), .Q(
        n2514) );
  AO22X1 U1633 ( .IN1(n3320), .IN2(n3621), .IN3(elem19[23]), .IN4(n3316), .Q(
        n2515) );
  AO22X1 U1634 ( .IN1(n3319), .IN2(n3624), .IN3(elem19[24]), .IN4(n3316), .Q(
        n2516) );
  AO22X1 U1635 ( .IN1(n3320), .IN2(n3627), .IN3(elem19[25]), .IN4(n3316), .Q(
        n2517) );
  AO22X1 U1636 ( .IN1(n3320), .IN2(n3630), .IN3(elem19[26]), .IN4(n3316), .Q(
        n2518) );
  AO22X1 U1637 ( .IN1(n3320), .IN2(n3633), .IN3(elem19[27]), .IN4(n3316), .Q(
        n2519) );
  AO22X1 U1638 ( .IN1(n3320), .IN2(n3636), .IN3(elem19[28]), .IN4(n3316), .Q(
        n2520) );
  AO22X1 U1639 ( .IN1(n3320), .IN2(n3639), .IN3(elem19[29]), .IN4(n3316), .Q(
        n2521) );
  AO22X1 U1640 ( .IN1(n3320), .IN2(n3642), .IN3(elem19[30]), .IN4(n3316), .Q(
        n2522) );
  AO22X1 U1641 ( .IN1(n3320), .IN2(n3645), .IN3(elem19[31]), .IN4(n3316), .Q(
        n2523) );
  AO22X1 U1642 ( .IN1(n3313), .IN2(n3553), .IN3(elem18[0]), .IN4(n2239), .Q(
        n2524) );
  AO22X1 U1643 ( .IN1(n3313), .IN2(n3556), .IN3(elem18[1]), .IN4(n2239), .Q(
        n2525) );
  AO22X1 U1644 ( .IN1(n3313), .IN2(n3559), .IN3(elem18[2]), .IN4(n2239), .Q(
        n2526) );
  AO22X1 U1645 ( .IN1(n3313), .IN2(n3562), .IN3(elem18[3]), .IN4(n2239), .Q(
        n2527) );
  AO22X1 U1646 ( .IN1(n3314), .IN2(n3565), .IN3(elem18[4]), .IN4(n2239), .Q(
        n2528) );
  AO22X1 U1647 ( .IN1(n3315), .IN2(n3568), .IN3(elem18[5]), .IN4(n2239), .Q(
        n2529) );
  AO22X1 U1648 ( .IN1(n3315), .IN2(n3571), .IN3(elem18[6]), .IN4(n2239), .Q(
        n2530) );
  AO22X1 U1649 ( .IN1(n3314), .IN2(n3574), .IN3(elem18[7]), .IN4(n2239), .Q(
        n2531) );
  AO22X1 U1650 ( .IN1(n3315), .IN2(n3577), .IN3(elem18[8]), .IN4(n3312), .Q(
        n2532) );
  AO22X1 U1651 ( .IN1(n3315), .IN2(n3580), .IN3(elem18[9]), .IN4(n3312), .Q(
        n2533) );
  AO22X1 U1652 ( .IN1(n3314), .IN2(n3583), .IN3(elem18[10]), .IN4(n3312), .Q(
        n2534) );
  AO22X1 U1653 ( .IN1(n3314), .IN2(n3586), .IN3(elem18[11]), .IN4(n3312), .Q(
        n2535) );
  AO22X1 U1654 ( .IN1(n3314), .IN2(n3588), .IN3(elem18[12]), .IN4(n3312), .Q(
        n2536) );
  AO22X1 U1655 ( .IN1(n3314), .IN2(n3591), .IN3(elem18[13]), .IN4(n3312), .Q(
        n2537) );
  AO22X1 U1656 ( .IN1(n3314), .IN2(n3594), .IN3(elem18[14]), .IN4(n3312), .Q(
        n2538) );
  AO22X1 U1657 ( .IN1(n3314), .IN2(n3597), .IN3(elem18[15]), .IN4(n3312), .Q(
        n2539) );
  AO22X1 U1658 ( .IN1(n3314), .IN2(n3600), .IN3(elem18[16]), .IN4(n3312), .Q(
        n2540) );
  AO22X1 U1659 ( .IN1(n3314), .IN2(n3603), .IN3(elem18[17]), .IN4(n3312), .Q(
        n2541) );
  AO22X1 U1660 ( .IN1(n3314), .IN2(n3606), .IN3(elem18[18]), .IN4(n3312), .Q(
        n2542) );
  AO22X1 U1661 ( .IN1(n3315), .IN2(n3609), .IN3(elem18[19]), .IN4(n3312), .Q(
        n2543) );
  AO22X1 U1662 ( .IN1(n3314), .IN2(n3612), .IN3(elem18[20]), .IN4(n3311), .Q(
        n2544) );
  AO22X1 U1663 ( .IN1(n3315), .IN2(n3615), .IN3(elem18[21]), .IN4(n3311), .Q(
        n2545) );
  AO22X1 U1664 ( .IN1(n3314), .IN2(n3618), .IN3(elem18[22]), .IN4(n3311), .Q(
        n2546) );
  AO22X1 U1665 ( .IN1(n3315), .IN2(n3621), .IN3(elem18[23]), .IN4(n3311), .Q(
        n2547) );
  AO22X1 U1666 ( .IN1(n3314), .IN2(n3624), .IN3(elem18[24]), .IN4(n3311), .Q(
        n2548) );
  AO22X1 U1667 ( .IN1(n3315), .IN2(n3627), .IN3(elem18[25]), .IN4(n3311), .Q(
        n2549) );
  AO22X1 U1668 ( .IN1(n3315), .IN2(n3630), .IN3(elem18[26]), .IN4(n3311), .Q(
        n2550) );
  AO22X1 U1669 ( .IN1(n3315), .IN2(n3633), .IN3(elem18[27]), .IN4(n3311), .Q(
        n2551) );
  AO22X1 U1670 ( .IN1(n3315), .IN2(n3636), .IN3(elem18[28]), .IN4(n3311), .Q(
        n2552) );
  AO22X1 U1671 ( .IN1(n3315), .IN2(n3639), .IN3(elem18[29]), .IN4(n3311), .Q(
        n2553) );
  AO22X1 U1672 ( .IN1(n3315), .IN2(n3642), .IN3(elem18[30]), .IN4(n3311), .Q(
        n2554) );
  AO22X1 U1673 ( .IN1(n3315), .IN2(n3645), .IN3(elem18[31]), .IN4(n3311), .Q(
        n2555) );
  AO22X1 U1674 ( .IN1(n3308), .IN2(n3553), .IN3(elem17[0]), .IN4(n2240), .Q(
        n2556) );
  AO22X1 U1675 ( .IN1(n3308), .IN2(n3556), .IN3(elem17[1]), .IN4(n2240), .Q(
        n2557) );
  AO22X1 U1676 ( .IN1(n3308), .IN2(n3559), .IN3(elem17[2]), .IN4(n2240), .Q(
        n2558) );
  AO22X1 U1677 ( .IN1(n3308), .IN2(n3562), .IN3(elem17[3]), .IN4(n2240), .Q(
        n2559) );
  AO22X1 U1678 ( .IN1(n3309), .IN2(n3565), .IN3(elem17[4]), .IN4(n2240), .Q(
        n2560) );
  AO22X1 U1679 ( .IN1(n3310), .IN2(n3568), .IN3(elem17[5]), .IN4(n2240), .Q(
        n2561) );
  AO22X1 U1680 ( .IN1(n3310), .IN2(n3571), .IN3(elem17[6]), .IN4(n2240), .Q(
        n2562) );
  AO22X1 U1681 ( .IN1(n3309), .IN2(n3574), .IN3(elem17[7]), .IN4(n2240), .Q(
        n2563) );
  AO22X1 U1682 ( .IN1(n3310), .IN2(n3577), .IN3(elem17[8]), .IN4(n3307), .Q(
        n2564) );
  AO22X1 U1683 ( .IN1(n3310), .IN2(n3580), .IN3(elem17[9]), .IN4(n3307), .Q(
        n2565) );
  AO22X1 U1684 ( .IN1(n3309), .IN2(n3583), .IN3(elem17[10]), .IN4(n3307), .Q(
        n2566) );
  AO22X1 U1685 ( .IN1(n3309), .IN2(n3586), .IN3(elem17[11]), .IN4(n3307), .Q(
        n2567) );
  AO22X1 U1686 ( .IN1(n3309), .IN2(n3588), .IN3(elem17[12]), .IN4(n3307), .Q(
        n2568) );
  AO22X1 U1687 ( .IN1(n3309), .IN2(n3591), .IN3(elem17[13]), .IN4(n3307), .Q(
        n2569) );
  AO22X1 U1688 ( .IN1(n3309), .IN2(n3594), .IN3(elem17[14]), .IN4(n3307), .Q(
        n2570) );
  AO22X1 U1689 ( .IN1(n3309), .IN2(n3597), .IN3(elem17[15]), .IN4(n3307), .Q(
        n2571) );
  AO22X1 U1690 ( .IN1(n3309), .IN2(n3600), .IN3(elem17[16]), .IN4(n3307), .Q(
        n2572) );
  AO22X1 U1691 ( .IN1(n3309), .IN2(n3603), .IN3(elem17[17]), .IN4(n3307), .Q(
        n2573) );
  AO22X1 U1692 ( .IN1(n3309), .IN2(n3606), .IN3(elem17[18]), .IN4(n3307), .Q(
        n2574) );
  AO22X1 U1693 ( .IN1(n3310), .IN2(n3609), .IN3(elem17[19]), .IN4(n3307), .Q(
        n2575) );
  AO22X1 U1694 ( .IN1(n3309), .IN2(n3612), .IN3(elem17[20]), .IN4(n3306), .Q(
        n2576) );
  AO22X1 U1695 ( .IN1(n3310), .IN2(n3615), .IN3(elem17[21]), .IN4(n3306), .Q(
        n2577) );
  AO22X1 U1696 ( .IN1(n3309), .IN2(n3618), .IN3(elem17[22]), .IN4(n3306), .Q(
        n2578) );
  AO22X1 U1697 ( .IN1(n3310), .IN2(n3621), .IN3(elem17[23]), .IN4(n3306), .Q(
        n2579) );
  AO22X1 U1698 ( .IN1(n3309), .IN2(n3624), .IN3(elem17[24]), .IN4(n3306), .Q(
        n2580) );
  AO22X1 U1699 ( .IN1(n3310), .IN2(n3627), .IN3(elem17[25]), .IN4(n3306), .Q(
        n2581) );
  AO22X1 U1700 ( .IN1(n3310), .IN2(n3630), .IN3(elem17[26]), .IN4(n3306), .Q(
        n2582) );
  AO22X1 U1701 ( .IN1(n3310), .IN2(n3633), .IN3(elem17[27]), .IN4(n3306), .Q(
        n2583) );
  AO22X1 U1702 ( .IN1(n3310), .IN2(n3636), .IN3(elem17[28]), .IN4(n3306), .Q(
        n2584) );
  AO22X1 U1703 ( .IN1(n3310), .IN2(n3639), .IN3(elem17[29]), .IN4(n3306), .Q(
        n2585) );
  AO22X1 U1704 ( .IN1(n3310), .IN2(n3642), .IN3(elem17[30]), .IN4(n3306), .Q(
        n2586) );
  AO22X1 U1705 ( .IN1(n3310), .IN2(n3645), .IN3(elem17[31]), .IN4(n3306), .Q(
        n2587) );
  AO22X1 U1706 ( .IN1(n3303), .IN2(n3553), .IN3(elem16[0]), .IN4(n2241), .Q(
        n2588) );
  AO22X1 U1707 ( .IN1(n3303), .IN2(n3556), .IN3(elem16[1]), .IN4(n2241), .Q(
        n2589) );
  AO22X1 U1708 ( .IN1(n3303), .IN2(n3559), .IN3(elem16[2]), .IN4(n2241), .Q(
        n2590) );
  AO22X1 U1709 ( .IN1(n3303), .IN2(n3562), .IN3(elem16[3]), .IN4(n2241), .Q(
        n2591) );
  AO22X1 U1710 ( .IN1(n3304), .IN2(n3565), .IN3(elem16[4]), .IN4(n2241), .Q(
        n2592) );
  AO22X1 U1711 ( .IN1(n3305), .IN2(n3568), .IN3(elem16[5]), .IN4(n2241), .Q(
        n2593) );
  AO22X1 U1712 ( .IN1(n3305), .IN2(n3571), .IN3(elem16[6]), .IN4(n2241), .Q(
        n2594) );
  AO22X1 U1713 ( .IN1(n3304), .IN2(n3574), .IN3(elem16[7]), .IN4(n2241), .Q(
        n2595) );
  AO22X1 U1714 ( .IN1(n3305), .IN2(n3577), .IN3(elem16[8]), .IN4(n3302), .Q(
        n2596) );
  AO22X1 U1715 ( .IN1(n3305), .IN2(n3580), .IN3(elem16[9]), .IN4(n3302), .Q(
        n2597) );
  AO22X1 U1716 ( .IN1(n3304), .IN2(n3583), .IN3(elem16[10]), .IN4(n3302), .Q(
        n2598) );
  AO22X1 U1717 ( .IN1(n3304), .IN2(n3586), .IN3(elem16[11]), .IN4(n3302), .Q(
        n2599) );
  AO22X1 U1718 ( .IN1(n3304), .IN2(n3589), .IN3(elem16[12]), .IN4(n3302), .Q(
        n2600) );
  AO22X1 U1719 ( .IN1(n3304), .IN2(n3592), .IN3(elem16[13]), .IN4(n3302), .Q(
        n2601) );
  AO22X1 U1720 ( .IN1(n3304), .IN2(n3595), .IN3(elem16[14]), .IN4(n3302), .Q(
        n2602) );
  AO22X1 U1721 ( .IN1(n3304), .IN2(n3598), .IN3(elem16[15]), .IN4(n3302), .Q(
        n2603) );
  AO22X1 U1722 ( .IN1(n3304), .IN2(n3601), .IN3(elem16[16]), .IN4(n3302), .Q(
        n2604) );
  AO22X1 U1723 ( .IN1(n3304), .IN2(n3604), .IN3(elem16[17]), .IN4(n3302), .Q(
        n2605) );
  AO22X1 U1724 ( .IN1(n3304), .IN2(n3607), .IN3(elem16[18]), .IN4(n3302), .Q(
        n2606) );
  AO22X1 U1725 ( .IN1(n3305), .IN2(n3610), .IN3(elem16[19]), .IN4(n3302), .Q(
        n2607) );
  AO22X1 U1726 ( .IN1(n3304), .IN2(n3613), .IN3(elem16[20]), .IN4(n3301), .Q(
        n2608) );
  AO22X1 U1727 ( .IN1(n3305), .IN2(n3616), .IN3(elem16[21]), .IN4(n3301), .Q(
        n2609) );
  AO22X1 U1728 ( .IN1(n3304), .IN2(n3619), .IN3(elem16[22]), .IN4(n3301), .Q(
        n2610) );
  AO22X1 U1729 ( .IN1(n3305), .IN2(n3622), .IN3(elem16[23]), .IN4(n3301), .Q(
        n2611) );
  AO22X1 U1730 ( .IN1(n3304), .IN2(n3625), .IN3(elem16[24]), .IN4(n3301), .Q(
        n2612) );
  AO22X1 U1731 ( .IN1(n3305), .IN2(n3628), .IN3(elem16[25]), .IN4(n3301), .Q(
        n2613) );
  AO22X1 U1732 ( .IN1(n3305), .IN2(n3631), .IN3(elem16[26]), .IN4(n3301), .Q(
        n2614) );
  AO22X1 U1733 ( .IN1(n3305), .IN2(n3634), .IN3(elem16[27]), .IN4(n3301), .Q(
        n2615) );
  AO22X1 U1734 ( .IN1(n3305), .IN2(n3637), .IN3(elem16[28]), .IN4(n3301), .Q(
        n2616) );
  AO22X1 U1735 ( .IN1(n3305), .IN2(n3640), .IN3(elem16[29]), .IN4(n3301), .Q(
        n2617) );
  AO22X1 U1736 ( .IN1(n3305), .IN2(n3643), .IN3(elem16[30]), .IN4(n3301), .Q(
        n2618) );
  AO22X1 U1737 ( .IN1(n3305), .IN2(n3646), .IN3(elem16[31]), .IN4(n3301), .Q(
        n2619) );
  AND2X1 U1738 ( .IN1(n2242), .IN2(n2230), .Q(n2238) );
  AO22X1 U1739 ( .IN1(n3298), .IN2(n3553), .IN3(elem15[0]), .IN4(n2243), .Q(
        n2620) );
  AO22X1 U1740 ( .IN1(n3298), .IN2(n3556), .IN3(elem15[1]), .IN4(n2243), .Q(
        n2621) );
  AO22X1 U1741 ( .IN1(n3298), .IN2(n3559), .IN3(elem15[2]), .IN4(n2243), .Q(
        n2622) );
  AO22X1 U1742 ( .IN1(n3298), .IN2(n3562), .IN3(elem15[3]), .IN4(n2243), .Q(
        n2623) );
  AO22X1 U1743 ( .IN1(n3299), .IN2(n3565), .IN3(elem15[4]), .IN4(n2243), .Q(
        n2624) );
  AO22X1 U1744 ( .IN1(n3300), .IN2(n3568), .IN3(elem15[5]), .IN4(n2243), .Q(
        n2625) );
  AO22X1 U1745 ( .IN1(n3300), .IN2(n3571), .IN3(elem15[6]), .IN4(n2243), .Q(
        n2626) );
  AO22X1 U1746 ( .IN1(n3299), .IN2(n3574), .IN3(elem15[7]), .IN4(n2243), .Q(
        n2627) );
  AO22X1 U1747 ( .IN1(n3300), .IN2(n3577), .IN3(elem15[8]), .IN4(n3297), .Q(
        n2628) );
  AO22X1 U1748 ( .IN1(n3300), .IN2(n3580), .IN3(elem15[9]), .IN4(n3297), .Q(
        n2629) );
  AO22X1 U1749 ( .IN1(n3299), .IN2(n3583), .IN3(elem15[10]), .IN4(n3297), .Q(
        n2630) );
  AO22X1 U1750 ( .IN1(n3299), .IN2(n3586), .IN3(elem15[11]), .IN4(n3297), .Q(
        n2631) );
  AO22X1 U1751 ( .IN1(n3299), .IN2(n3589), .IN3(elem15[12]), .IN4(n3297), .Q(
        n2632) );
  AO22X1 U1752 ( .IN1(n3299), .IN2(n3592), .IN3(elem15[13]), .IN4(n3297), .Q(
        n2633) );
  AO22X1 U1753 ( .IN1(n3299), .IN2(n3595), .IN3(elem15[14]), .IN4(n3297), .Q(
        n2634) );
  AO22X1 U1754 ( .IN1(n3299), .IN2(n3598), .IN3(elem15[15]), .IN4(n3297), .Q(
        n2635) );
  AO22X1 U1755 ( .IN1(n3299), .IN2(n3601), .IN3(elem15[16]), .IN4(n3297), .Q(
        n2636) );
  AO22X1 U1756 ( .IN1(n3299), .IN2(n3604), .IN3(elem15[17]), .IN4(n3297), .Q(
        n2637) );
  AO22X1 U1757 ( .IN1(n3299), .IN2(n3607), .IN3(elem15[18]), .IN4(n3297), .Q(
        n2638) );
  AO22X1 U1758 ( .IN1(n3300), .IN2(n3610), .IN3(elem15[19]), .IN4(n3297), .Q(
        n2639) );
  AO22X1 U1759 ( .IN1(n3299), .IN2(n3613), .IN3(elem15[20]), .IN4(n3296), .Q(
        n2640) );
  AO22X1 U1760 ( .IN1(n3300), .IN2(n3616), .IN3(elem15[21]), .IN4(n3296), .Q(
        n2641) );
  AO22X1 U1761 ( .IN1(n3299), .IN2(n3619), .IN3(elem15[22]), .IN4(n3296), .Q(
        n2642) );
  AO22X1 U1762 ( .IN1(n3300), .IN2(n3622), .IN3(elem15[23]), .IN4(n3296), .Q(
        n2643) );
  AO22X1 U1763 ( .IN1(n3299), .IN2(n3625), .IN3(elem15[24]), .IN4(n3296), .Q(
        n2644) );
  AO22X1 U1764 ( .IN1(n3300), .IN2(n3628), .IN3(elem15[25]), .IN4(n3296), .Q(
        n2645) );
  AO22X1 U1765 ( .IN1(n3300), .IN2(n3631), .IN3(elem15[26]), .IN4(n3296), .Q(
        n2646) );
  AO22X1 U1766 ( .IN1(n3300), .IN2(n3634), .IN3(elem15[27]), .IN4(n3296), .Q(
        n2647) );
  AO22X1 U1767 ( .IN1(n3300), .IN2(n3637), .IN3(elem15[28]), .IN4(n3296), .Q(
        n2648) );
  AO22X1 U1768 ( .IN1(n3300), .IN2(n3640), .IN3(elem15[29]), .IN4(n3296), .Q(
        n2649) );
  AO22X1 U1769 ( .IN1(n3300), .IN2(n3643), .IN3(elem15[30]), .IN4(n3296), .Q(
        n2650) );
  AO22X1 U1770 ( .IN1(n3300), .IN2(n3646), .IN3(elem15[31]), .IN4(n3296), .Q(
        n2651) );
  AO22X1 U1771 ( .IN1(n3293), .IN2(n3553), .IN3(elem14[0]), .IN4(n2245), .Q(
        n2652) );
  AO22X1 U1772 ( .IN1(n3293), .IN2(n3556), .IN3(elem14[1]), .IN4(n2245), .Q(
        n2653) );
  AO22X1 U1773 ( .IN1(n3293), .IN2(n3559), .IN3(elem14[2]), .IN4(n2245), .Q(
        n2654) );
  AO22X1 U1774 ( .IN1(n3293), .IN2(n3562), .IN3(elem14[3]), .IN4(n2245), .Q(
        n2655) );
  AO22X1 U1775 ( .IN1(n3294), .IN2(n3565), .IN3(elem14[4]), .IN4(n2245), .Q(
        n2656) );
  AO22X1 U1776 ( .IN1(n3295), .IN2(n3568), .IN3(elem14[5]), .IN4(n2245), .Q(
        n2657) );
  AO22X1 U1777 ( .IN1(n3295), .IN2(n3571), .IN3(elem14[6]), .IN4(n2245), .Q(
        n2658) );
  AO22X1 U1778 ( .IN1(n3294), .IN2(n3574), .IN3(elem14[7]), .IN4(n2245), .Q(
        n2659) );
  AO22X1 U1779 ( .IN1(n3295), .IN2(n3577), .IN3(elem14[8]), .IN4(n3292), .Q(
        n2660) );
  AO22X1 U1780 ( .IN1(n3295), .IN2(n3580), .IN3(elem14[9]), .IN4(n3292), .Q(
        n2661) );
  AO22X1 U1781 ( .IN1(n3294), .IN2(n3583), .IN3(elem14[10]), .IN4(n3292), .Q(
        n2662) );
  AO22X1 U1782 ( .IN1(n3294), .IN2(n3586), .IN3(elem14[11]), .IN4(n3292), .Q(
        n2663) );
  AO22X1 U1783 ( .IN1(n3294), .IN2(n3589), .IN3(elem14[12]), .IN4(n3292), .Q(
        n2664) );
  AO22X1 U1784 ( .IN1(n3294), .IN2(n3592), .IN3(elem14[13]), .IN4(n3292), .Q(
        n2665) );
  AO22X1 U1785 ( .IN1(n3294), .IN2(n3595), .IN3(elem14[14]), .IN4(n3292), .Q(
        n2666) );
  AO22X1 U1786 ( .IN1(n3294), .IN2(n3598), .IN3(elem14[15]), .IN4(n3292), .Q(
        n2667) );
  AO22X1 U1787 ( .IN1(n3294), .IN2(n3601), .IN3(elem14[16]), .IN4(n3292), .Q(
        n2668) );
  AO22X1 U1788 ( .IN1(n3294), .IN2(n3604), .IN3(elem14[17]), .IN4(n3292), .Q(
        n2669) );
  AO22X1 U1789 ( .IN1(n3294), .IN2(n3607), .IN3(elem14[18]), .IN4(n3292), .Q(
        n2670) );
  AO22X1 U1790 ( .IN1(n3295), .IN2(n3610), .IN3(elem14[19]), .IN4(n3292), .Q(
        n2671) );
  AO22X1 U1791 ( .IN1(n3294), .IN2(n3613), .IN3(elem14[20]), .IN4(n3291), .Q(
        n2672) );
  AO22X1 U1792 ( .IN1(n3295), .IN2(n3616), .IN3(elem14[21]), .IN4(n3291), .Q(
        n2673) );
  AO22X1 U1793 ( .IN1(n3294), .IN2(n3619), .IN3(elem14[22]), .IN4(n3291), .Q(
        n2674) );
  AO22X1 U1794 ( .IN1(n3295), .IN2(n3622), .IN3(elem14[23]), .IN4(n3291), .Q(
        n2675) );
  AO22X1 U1795 ( .IN1(n3294), .IN2(n3625), .IN3(elem14[24]), .IN4(n3291), .Q(
        n2676) );
  AO22X1 U1796 ( .IN1(n3295), .IN2(n3628), .IN3(elem14[25]), .IN4(n3291), .Q(
        n2677) );
  AO22X1 U1797 ( .IN1(n3295), .IN2(n3631), .IN3(elem14[26]), .IN4(n3291), .Q(
        n2678) );
  AO22X1 U1798 ( .IN1(n3295), .IN2(n3634), .IN3(elem14[27]), .IN4(n3291), .Q(
        n2679) );
  AO22X1 U1799 ( .IN1(n3295), .IN2(n3637), .IN3(elem14[28]), .IN4(n3291), .Q(
        n2680) );
  AO22X1 U1800 ( .IN1(n3295), .IN2(n3640), .IN3(elem14[29]), .IN4(n3291), .Q(
        n2681) );
  AO22X1 U1801 ( .IN1(n3295), .IN2(n3643), .IN3(elem14[30]), .IN4(n3291), .Q(
        n2682) );
  AO22X1 U1802 ( .IN1(n3295), .IN2(n3646), .IN3(elem14[31]), .IN4(n3291), .Q(
        n2683) );
  AO22X1 U1803 ( .IN1(n3288), .IN2(n3553), .IN3(elem13[0]), .IN4(n2246), .Q(
        n2684) );
  AO22X1 U1804 ( .IN1(n3288), .IN2(n3556), .IN3(elem13[1]), .IN4(n2246), .Q(
        n2685) );
  AO22X1 U1805 ( .IN1(n3288), .IN2(n3559), .IN3(elem13[2]), .IN4(n2246), .Q(
        n2686) );
  AO22X1 U1806 ( .IN1(n3288), .IN2(n3562), .IN3(elem13[3]), .IN4(n2246), .Q(
        n2687) );
  AO22X1 U1807 ( .IN1(n3289), .IN2(n3565), .IN3(elem13[4]), .IN4(n2246), .Q(
        n2688) );
  AO22X1 U1808 ( .IN1(n3290), .IN2(n3568), .IN3(elem13[5]), .IN4(n2246), .Q(
        n2689) );
  AO22X1 U1809 ( .IN1(n3290), .IN2(n3571), .IN3(elem13[6]), .IN4(n2246), .Q(
        n2690) );
  AO22X1 U1810 ( .IN1(n3289), .IN2(n3574), .IN3(elem13[7]), .IN4(n2246), .Q(
        n2691) );
  AO22X1 U1811 ( .IN1(n3290), .IN2(n3577), .IN3(elem13[8]), .IN4(n3287), .Q(
        n2692) );
  AO22X1 U1812 ( .IN1(n3290), .IN2(n3580), .IN3(elem13[9]), .IN4(n3287), .Q(
        n2693) );
  AO22X1 U1813 ( .IN1(n3289), .IN2(n3583), .IN3(elem13[10]), .IN4(n3287), .Q(
        n2694) );
  AO22X1 U1814 ( .IN1(n3289), .IN2(n3586), .IN3(elem13[11]), .IN4(n3287), .Q(
        n2695) );
  AO22X1 U1815 ( .IN1(n3289), .IN2(n3589), .IN3(elem13[12]), .IN4(n3287), .Q(
        n2696) );
  AO22X1 U1816 ( .IN1(n3289), .IN2(n3592), .IN3(elem13[13]), .IN4(n3287), .Q(
        n2697) );
  AO22X1 U1817 ( .IN1(n3289), .IN2(n3595), .IN3(elem13[14]), .IN4(n3287), .Q(
        n2698) );
  AO22X1 U1818 ( .IN1(n3289), .IN2(n3598), .IN3(elem13[15]), .IN4(n3287), .Q(
        n2699) );
  AO22X1 U1819 ( .IN1(n3289), .IN2(n3601), .IN3(elem13[16]), .IN4(n3287), .Q(
        n2700) );
  AO22X1 U1820 ( .IN1(n3289), .IN2(n3604), .IN3(elem13[17]), .IN4(n3287), .Q(
        n2701) );
  AO22X1 U1821 ( .IN1(n3289), .IN2(n3607), .IN3(elem13[18]), .IN4(n3287), .Q(
        n2702) );
  AO22X1 U1822 ( .IN1(n3290), .IN2(n3610), .IN3(elem13[19]), .IN4(n3287), .Q(
        n2703) );
  AO22X1 U1823 ( .IN1(n3289), .IN2(n3613), .IN3(elem13[20]), .IN4(n3286), .Q(
        n2704) );
  AO22X1 U1824 ( .IN1(n3290), .IN2(n3616), .IN3(elem13[21]), .IN4(n3286), .Q(
        n2705) );
  AO22X1 U1825 ( .IN1(n3289), .IN2(n3619), .IN3(elem13[22]), .IN4(n3286), .Q(
        n2706) );
  AO22X1 U1826 ( .IN1(n3290), .IN2(n3622), .IN3(elem13[23]), .IN4(n3286), .Q(
        n2707) );
  AO22X1 U1827 ( .IN1(n3289), .IN2(n3625), .IN3(elem13[24]), .IN4(n3286), .Q(
        n2708) );
  AO22X1 U1828 ( .IN1(n3290), .IN2(n3628), .IN3(elem13[25]), .IN4(n3286), .Q(
        n2709) );
  AO22X1 U1829 ( .IN1(n3290), .IN2(n3631), .IN3(elem13[26]), .IN4(n3286), .Q(
        n2710) );
  AO22X1 U1830 ( .IN1(n3290), .IN2(n3634), .IN3(elem13[27]), .IN4(n3286), .Q(
        n2711) );
  AO22X1 U1831 ( .IN1(n3290), .IN2(n3637), .IN3(elem13[28]), .IN4(n3286), .Q(
        n2712) );
  AO22X1 U1832 ( .IN1(n3290), .IN2(n3640), .IN3(elem13[29]), .IN4(n3286), .Q(
        n2713) );
  AO22X1 U1833 ( .IN1(n3290), .IN2(n3643), .IN3(elem13[30]), .IN4(n3286), .Q(
        n2714) );
  AO22X1 U1834 ( .IN1(n3290), .IN2(n3646), .IN3(elem13[31]), .IN4(n3286), .Q(
        n2715) );
  AO22X1 U1835 ( .IN1(n3283), .IN2(n3553), .IN3(elem12[0]), .IN4(n2247), .Q(
        n2716) );
  AO22X1 U1836 ( .IN1(n3283), .IN2(n3556), .IN3(elem12[1]), .IN4(n2247), .Q(
        n2717) );
  AO22X1 U1837 ( .IN1(n3283), .IN2(n3559), .IN3(elem12[2]), .IN4(n2247), .Q(
        n2718) );
  AO22X1 U1838 ( .IN1(n3283), .IN2(n3562), .IN3(elem12[3]), .IN4(n2247), .Q(
        n2719) );
  AO22X1 U1839 ( .IN1(n3284), .IN2(n3565), .IN3(elem12[4]), .IN4(n2247), .Q(
        n2720) );
  AO22X1 U1840 ( .IN1(n3285), .IN2(n3568), .IN3(elem12[5]), .IN4(n2247), .Q(
        n2721) );
  AO22X1 U1841 ( .IN1(n3285), .IN2(n3571), .IN3(elem12[6]), .IN4(n2247), .Q(
        n2722) );
  AO22X1 U1842 ( .IN1(n3284), .IN2(n3574), .IN3(elem12[7]), .IN4(n2247), .Q(
        n2723) );
  AO22X1 U1843 ( .IN1(n3285), .IN2(n3577), .IN3(elem12[8]), .IN4(n3282), .Q(
        n2724) );
  AO22X1 U1844 ( .IN1(n3285), .IN2(n3580), .IN3(elem12[9]), .IN4(n3282), .Q(
        n2725) );
  AO22X1 U1845 ( .IN1(n3284), .IN2(n3583), .IN3(elem12[10]), .IN4(n3282), .Q(
        n2726) );
  AO22X1 U1846 ( .IN1(n3284), .IN2(n3586), .IN3(elem12[11]), .IN4(n3282), .Q(
        n2727) );
  AO22X1 U1847 ( .IN1(n3284), .IN2(n3589), .IN3(elem12[12]), .IN4(n3282), .Q(
        n2728) );
  AO22X1 U1848 ( .IN1(n3284), .IN2(n3592), .IN3(elem12[13]), .IN4(n3282), .Q(
        n2729) );
  AO22X1 U1849 ( .IN1(n3284), .IN2(n3595), .IN3(elem12[14]), .IN4(n3282), .Q(
        n2730) );
  AO22X1 U1850 ( .IN1(n3284), .IN2(n3598), .IN3(elem12[15]), .IN4(n3282), .Q(
        n2731) );
  AO22X1 U1851 ( .IN1(n3284), .IN2(n3601), .IN3(elem12[16]), .IN4(n3282), .Q(
        n2732) );
  AO22X1 U1852 ( .IN1(n3284), .IN2(n3604), .IN3(elem12[17]), .IN4(n3282), .Q(
        n2733) );
  AO22X1 U1853 ( .IN1(n3284), .IN2(n3607), .IN3(elem12[18]), .IN4(n3282), .Q(
        n2734) );
  AO22X1 U1854 ( .IN1(n3285), .IN2(n3610), .IN3(elem12[19]), .IN4(n3282), .Q(
        n2735) );
  AO22X1 U1855 ( .IN1(n3284), .IN2(n3613), .IN3(elem12[20]), .IN4(n3281), .Q(
        n2736) );
  AO22X1 U1856 ( .IN1(n3285), .IN2(n3616), .IN3(elem12[21]), .IN4(n3281), .Q(
        n2737) );
  AO22X1 U1857 ( .IN1(n3284), .IN2(n3619), .IN3(elem12[22]), .IN4(n3281), .Q(
        n2738) );
  AO22X1 U1858 ( .IN1(n3285), .IN2(n3622), .IN3(elem12[23]), .IN4(n3281), .Q(
        n2739) );
  AO22X1 U1859 ( .IN1(n3284), .IN2(n3625), .IN3(elem12[24]), .IN4(n3281), .Q(
        n2740) );
  AO22X1 U1860 ( .IN1(n3285), .IN2(n3628), .IN3(elem12[25]), .IN4(n3281), .Q(
        n2741) );
  AO22X1 U1861 ( .IN1(n3285), .IN2(n3631), .IN3(elem12[26]), .IN4(n3281), .Q(
        n2742) );
  AO22X1 U1862 ( .IN1(n3285), .IN2(n3634), .IN3(elem12[27]), .IN4(n3281), .Q(
        n2743) );
  AO22X1 U1863 ( .IN1(n3285), .IN2(n3637), .IN3(elem12[28]), .IN4(n3281), .Q(
        n2744) );
  AO22X1 U1864 ( .IN1(n3285), .IN2(n3640), .IN3(elem12[29]), .IN4(n3281), .Q(
        n2745) );
  AO22X1 U1865 ( .IN1(n3285), .IN2(n3643), .IN3(elem12[30]), .IN4(n3281), .Q(
        n2746) );
  AO22X1 U1866 ( .IN1(n3285), .IN2(n3646), .IN3(elem12[31]), .IN4(n3281), .Q(
        n2747) );
  AND2X1 U1867 ( .IN1(n2248), .IN2(n2249), .Q(n2244) );
  AO22X1 U1868 ( .IN1(n3278), .IN2(n3553), .IN3(elem11[0]), .IN4(n2250), .Q(
        n2748) );
  AO22X1 U1869 ( .IN1(n3278), .IN2(n3556), .IN3(elem11[1]), .IN4(n2250), .Q(
        n2749) );
  AO22X1 U1870 ( .IN1(n3278), .IN2(n3559), .IN3(elem11[2]), .IN4(n2250), .Q(
        n2750) );
  AO22X1 U1871 ( .IN1(n3278), .IN2(n3562), .IN3(elem11[3]), .IN4(n2250), .Q(
        n2751) );
  AO22X1 U1872 ( .IN1(n3279), .IN2(n3565), .IN3(elem11[4]), .IN4(n2250), .Q(
        n2752) );
  AO22X1 U1873 ( .IN1(n3280), .IN2(n3568), .IN3(elem11[5]), .IN4(n2250), .Q(
        n2753) );
  AO22X1 U1874 ( .IN1(n3280), .IN2(n3571), .IN3(elem11[6]), .IN4(n2250), .Q(
        n2754) );
  AO22X1 U1875 ( .IN1(n3279), .IN2(n3574), .IN3(elem11[7]), .IN4(n2250), .Q(
        n2755) );
  AO22X1 U1876 ( .IN1(n3280), .IN2(n3577), .IN3(elem11[8]), .IN4(n3277), .Q(
        n2756) );
  AO22X1 U1877 ( .IN1(n3280), .IN2(n3580), .IN3(elem11[9]), .IN4(n3277), .Q(
        n2757) );
  AO22X1 U1878 ( .IN1(n3279), .IN2(n3583), .IN3(elem11[10]), .IN4(n3277), .Q(
        n2758) );
  AO22X1 U1879 ( .IN1(n3279), .IN2(n3586), .IN3(elem11[11]), .IN4(n3277), .Q(
        n2759) );
  AO22X1 U1880 ( .IN1(n3279), .IN2(n3589), .IN3(elem11[12]), .IN4(n3277), .Q(
        n2760) );
  AO22X1 U1881 ( .IN1(n3279), .IN2(n3592), .IN3(elem11[13]), .IN4(n3277), .Q(
        n2761) );
  AO22X1 U1882 ( .IN1(n3279), .IN2(n3595), .IN3(elem11[14]), .IN4(n3277), .Q(
        n2762) );
  AO22X1 U1883 ( .IN1(n3279), .IN2(n3598), .IN3(elem11[15]), .IN4(n3277), .Q(
        n2763) );
  AO22X1 U1884 ( .IN1(n3279), .IN2(n3601), .IN3(elem11[16]), .IN4(n3277), .Q(
        n2764) );
  AO22X1 U1885 ( .IN1(n3279), .IN2(n3604), .IN3(elem11[17]), .IN4(n3277), .Q(
        n2765) );
  AO22X1 U1886 ( .IN1(n3279), .IN2(n3607), .IN3(elem11[18]), .IN4(n3277), .Q(
        n2766) );
  AO22X1 U1887 ( .IN1(n3280), .IN2(n3610), .IN3(elem11[19]), .IN4(n3277), .Q(
        n2767) );
  AO22X1 U1888 ( .IN1(n3279), .IN2(n3613), .IN3(elem11[20]), .IN4(n3276), .Q(
        n2768) );
  AO22X1 U1889 ( .IN1(n3280), .IN2(n3616), .IN3(elem11[21]), .IN4(n3276), .Q(
        n2769) );
  AO22X1 U1890 ( .IN1(n3279), .IN2(n3619), .IN3(elem11[22]), .IN4(n3276), .Q(
        n2770) );
  AO22X1 U1891 ( .IN1(n3280), .IN2(n3622), .IN3(elem11[23]), .IN4(n3276), .Q(
        n2771) );
  AO22X1 U1892 ( .IN1(n3279), .IN2(n3625), .IN3(elem11[24]), .IN4(n3276), .Q(
        n2772) );
  AO22X1 U1893 ( .IN1(n3280), .IN2(n3628), .IN3(elem11[25]), .IN4(n3276), .Q(
        n2773) );
  AO22X1 U1894 ( .IN1(n3280), .IN2(n3631), .IN3(elem11[26]), .IN4(n3276), .Q(
        n2774) );
  AO22X1 U1895 ( .IN1(n3280), .IN2(n3634), .IN3(elem11[27]), .IN4(n3276), .Q(
        n2775) );
  AO22X1 U1896 ( .IN1(n3280), .IN2(n3637), .IN3(elem11[28]), .IN4(n3276), .Q(
        n2776) );
  AO22X1 U1897 ( .IN1(n3280), .IN2(n3640), .IN3(elem11[29]), .IN4(n3276), .Q(
        n2777) );
  AO22X1 U1898 ( .IN1(n3280), .IN2(n3643), .IN3(elem11[30]), .IN4(n3276), .Q(
        n2778) );
  AO22X1 U1899 ( .IN1(n3280), .IN2(n3646), .IN3(elem11[31]), .IN4(n3276), .Q(
        n2779) );
  AO22X1 U1900 ( .IN1(n3273), .IN2(n3553), .IN3(elem10[0]), .IN4(n2252), .Q(
        n2780) );
  AO22X1 U1901 ( .IN1(n3273), .IN2(n3556), .IN3(elem10[1]), .IN4(n2252), .Q(
        n2781) );
  AO22X1 U1902 ( .IN1(n3273), .IN2(n3559), .IN3(elem10[2]), .IN4(n2252), .Q(
        n2782) );
  AO22X1 U1903 ( .IN1(n3273), .IN2(n3562), .IN3(elem10[3]), .IN4(n2252), .Q(
        n2783) );
  AO22X1 U1904 ( .IN1(n3274), .IN2(n3565), .IN3(elem10[4]), .IN4(n2252), .Q(
        n2784) );
  AO22X1 U1905 ( .IN1(n3275), .IN2(n3568), .IN3(elem10[5]), .IN4(n2252), .Q(
        n2785) );
  AO22X1 U1906 ( .IN1(n3275), .IN2(n3571), .IN3(elem10[6]), .IN4(n2252), .Q(
        n2786) );
  AO22X1 U1907 ( .IN1(n3274), .IN2(n3574), .IN3(elem10[7]), .IN4(n2252), .Q(
        n2787) );
  AO22X1 U1908 ( .IN1(n3275), .IN2(n3577), .IN3(elem10[8]), .IN4(n3272), .Q(
        n2788) );
  AO22X1 U1909 ( .IN1(n3275), .IN2(n3580), .IN3(elem10[9]), .IN4(n3272), .Q(
        n2789) );
  AO22X1 U1910 ( .IN1(n3274), .IN2(n3583), .IN3(elem10[10]), .IN4(n3272), .Q(
        n2790) );
  AO22X1 U1911 ( .IN1(n3274), .IN2(n3586), .IN3(elem10[11]), .IN4(n3272), .Q(
        n2791) );
  AO22X1 U1912 ( .IN1(n3274), .IN2(n3589), .IN3(elem10[12]), .IN4(n3272), .Q(
        n2792) );
  AO22X1 U1913 ( .IN1(n3274), .IN2(n3592), .IN3(elem10[13]), .IN4(n3272), .Q(
        n2793) );
  AO22X1 U1914 ( .IN1(n3274), .IN2(n3595), .IN3(elem10[14]), .IN4(n3272), .Q(
        n2794) );
  AO22X1 U1915 ( .IN1(n3274), .IN2(n3598), .IN3(elem10[15]), .IN4(n3272), .Q(
        n2795) );
  AO22X1 U1916 ( .IN1(n3274), .IN2(n3601), .IN3(elem10[16]), .IN4(n3272), .Q(
        n2796) );
  AO22X1 U1917 ( .IN1(n3274), .IN2(n3604), .IN3(elem10[17]), .IN4(n3272), .Q(
        n2797) );
  AO22X1 U1918 ( .IN1(n3274), .IN2(n3607), .IN3(elem10[18]), .IN4(n3272), .Q(
        n2798) );
  AO22X1 U1919 ( .IN1(n3275), .IN2(n3610), .IN3(elem10[19]), .IN4(n3272), .Q(
        n2799) );
  AO22X1 U1920 ( .IN1(n3274), .IN2(n3613), .IN3(elem10[20]), .IN4(n3271), .Q(
        n2800) );
  AO22X1 U1921 ( .IN1(n3275), .IN2(n3616), .IN3(elem10[21]), .IN4(n3271), .Q(
        n2801) );
  AO22X1 U1922 ( .IN1(n3274), .IN2(n3619), .IN3(elem10[22]), .IN4(n3271), .Q(
        n2802) );
  AO22X1 U1923 ( .IN1(n3275), .IN2(n3622), .IN3(elem10[23]), .IN4(n3271), .Q(
        n2803) );
  AO22X1 U1924 ( .IN1(n3274), .IN2(n3625), .IN3(elem10[24]), .IN4(n3271), .Q(
        n2804) );
  AO22X1 U1925 ( .IN1(n3275), .IN2(n3628), .IN3(elem10[25]), .IN4(n3271), .Q(
        n2805) );
  AO22X1 U1926 ( .IN1(n3275), .IN2(n3631), .IN3(elem10[26]), .IN4(n3271), .Q(
        n2806) );
  AO22X1 U1927 ( .IN1(n3275), .IN2(n3634), .IN3(elem10[27]), .IN4(n3271), .Q(
        n2807) );
  AO22X1 U1928 ( .IN1(n3275), .IN2(n3637), .IN3(elem10[28]), .IN4(n3271), .Q(
        n2808) );
  AO22X1 U1929 ( .IN1(n3275), .IN2(n3640), .IN3(elem10[29]), .IN4(n3271), .Q(
        n2809) );
  AO22X1 U1930 ( .IN1(n3275), .IN2(n3643), .IN3(elem10[30]), .IN4(n3271), .Q(
        n2810) );
  AO22X1 U1931 ( .IN1(n3275), .IN2(n3646), .IN3(elem10[31]), .IN4(n3271), .Q(
        n2811) );
  AO22X1 U1932 ( .IN1(n3268), .IN2(n3553), .IN3(elem09[0]), .IN4(n2253), .Q(
        n2812) );
  AO22X1 U1933 ( .IN1(n3268), .IN2(n3556), .IN3(elem09[1]), .IN4(n2253), .Q(
        n2813) );
  AO22X1 U1934 ( .IN1(n3268), .IN2(n3559), .IN3(elem09[2]), .IN4(n2253), .Q(
        n2814) );
  AO22X1 U1935 ( .IN1(n3268), .IN2(n3562), .IN3(elem09[3]), .IN4(n2253), .Q(
        n2815) );
  AO22X1 U1936 ( .IN1(n3269), .IN2(n3565), .IN3(elem09[4]), .IN4(n2253), .Q(
        n2816) );
  AO22X1 U1937 ( .IN1(n3270), .IN2(n3568), .IN3(elem09[5]), .IN4(n2253), .Q(
        n2817) );
  AO22X1 U1938 ( .IN1(n3270), .IN2(n3571), .IN3(elem09[6]), .IN4(n2253), .Q(
        n2818) );
  AO22X1 U1939 ( .IN1(n3269), .IN2(n3574), .IN3(elem09[7]), .IN4(n2253), .Q(
        n2819) );
  AO22X1 U1940 ( .IN1(n3270), .IN2(n3577), .IN3(elem09[8]), .IN4(n3267), .Q(
        n2820) );
  AO22X1 U1941 ( .IN1(n3270), .IN2(n3580), .IN3(elem09[9]), .IN4(n3267), .Q(
        n2821) );
  AO22X1 U1942 ( .IN1(n3269), .IN2(n3583), .IN3(elem09[10]), .IN4(n3267), .Q(
        n2822) );
  AO22X1 U1943 ( .IN1(n3269), .IN2(n3586), .IN3(elem09[11]), .IN4(n3267), .Q(
        n2823) );
  AO22X1 U1944 ( .IN1(n3269), .IN2(n3589), .IN3(elem09[12]), .IN4(n3267), .Q(
        n2824) );
  AO22X1 U1945 ( .IN1(n3269), .IN2(n3592), .IN3(elem09[13]), .IN4(n3267), .Q(
        n2825) );
  AO22X1 U1946 ( .IN1(n3269), .IN2(n3595), .IN3(elem09[14]), .IN4(n3267), .Q(
        n2826) );
  AO22X1 U1947 ( .IN1(n3269), .IN2(n3598), .IN3(elem09[15]), .IN4(n3267), .Q(
        n2827) );
  AO22X1 U1948 ( .IN1(n3269), .IN2(n3601), .IN3(elem09[16]), .IN4(n3267), .Q(
        n2828) );
  AO22X1 U1949 ( .IN1(n3269), .IN2(n3604), .IN3(elem09[17]), .IN4(n3267), .Q(
        n2829) );
  AO22X1 U1950 ( .IN1(n3269), .IN2(n3607), .IN3(elem09[18]), .IN4(n3267), .Q(
        n2830) );
  AO22X1 U1951 ( .IN1(n3270), .IN2(n3610), .IN3(elem09[19]), .IN4(n3267), .Q(
        n2831) );
  AO22X1 U1952 ( .IN1(n3269), .IN2(n3613), .IN3(elem09[20]), .IN4(n3266), .Q(
        n2832) );
  AO22X1 U1953 ( .IN1(n3270), .IN2(n3616), .IN3(elem09[21]), .IN4(n3266), .Q(
        n2833) );
  AO22X1 U1954 ( .IN1(n3269), .IN2(n3619), .IN3(elem09[22]), .IN4(n3266), .Q(
        n2834) );
  AO22X1 U1955 ( .IN1(n3270), .IN2(n3622), .IN3(elem09[23]), .IN4(n3266), .Q(
        n2835) );
  AO22X1 U1956 ( .IN1(n3269), .IN2(n3625), .IN3(elem09[24]), .IN4(n3266), .Q(
        n2836) );
  AO22X1 U1957 ( .IN1(n3270), .IN2(n3628), .IN3(elem09[25]), .IN4(n3266), .Q(
        n2837) );
  AO22X1 U1958 ( .IN1(n3270), .IN2(n3631), .IN3(elem09[26]), .IN4(n3266), .Q(
        n2838) );
  AO22X1 U1959 ( .IN1(n3270), .IN2(n3634), .IN3(elem09[27]), .IN4(n3266), .Q(
        n2839) );
  AO22X1 U1960 ( .IN1(n3270), .IN2(n3637), .IN3(elem09[28]), .IN4(n3266), .Q(
        n2840) );
  AO22X1 U1961 ( .IN1(n3270), .IN2(n3640), .IN3(elem09[29]), .IN4(n3266), .Q(
        n2841) );
  AO22X1 U1962 ( .IN1(n3270), .IN2(n3643), .IN3(elem09[30]), .IN4(n3266), .Q(
        n2842) );
  AO22X1 U1963 ( .IN1(n3270), .IN2(n3646), .IN3(elem09[31]), .IN4(n3266), .Q(
        n2843) );
  AO22X1 U1964 ( .IN1(n3263), .IN2(n3553), .IN3(elem08[0]), .IN4(n2254), .Q(
        n2844) );
  AO22X1 U1965 ( .IN1(n3263), .IN2(n3556), .IN3(elem08[1]), .IN4(n2254), .Q(
        n2845) );
  AO22X1 U1966 ( .IN1(n3263), .IN2(n3559), .IN3(elem08[2]), .IN4(n2254), .Q(
        n2846) );
  AO22X1 U1967 ( .IN1(n3263), .IN2(n3562), .IN3(elem08[3]), .IN4(n2254), .Q(
        n2847) );
  AO22X1 U1968 ( .IN1(n3264), .IN2(n3565), .IN3(elem08[4]), .IN4(n2254), .Q(
        n2848) );
  AO22X1 U1969 ( .IN1(n3265), .IN2(n3568), .IN3(elem08[5]), .IN4(n2254), .Q(
        n2849) );
  AO22X1 U1970 ( .IN1(n3265), .IN2(n3571), .IN3(elem08[6]), .IN4(n2254), .Q(
        n2850) );
  AO22X1 U1971 ( .IN1(n3264), .IN2(n3574), .IN3(elem08[7]), .IN4(n2254), .Q(
        n2851) );
  AO22X1 U1972 ( .IN1(n3265), .IN2(n3577), .IN3(elem08[8]), .IN4(n3262), .Q(
        n2852) );
  AO22X1 U1973 ( .IN1(n3265), .IN2(n3580), .IN3(elem08[9]), .IN4(n3262), .Q(
        n2853) );
  AO22X1 U1974 ( .IN1(n3264), .IN2(n3583), .IN3(elem08[10]), .IN4(n3262), .Q(
        n2854) );
  AO22X1 U1975 ( .IN1(n3264), .IN2(n3586), .IN3(elem08[11]), .IN4(n3262), .Q(
        n2855) );
  AO22X1 U1976 ( .IN1(n3264), .IN2(n3589), .IN3(elem08[12]), .IN4(n3262), .Q(
        n2856) );
  AO22X1 U1977 ( .IN1(n3264), .IN2(n3592), .IN3(elem08[13]), .IN4(n3262), .Q(
        n2857) );
  AO22X1 U1978 ( .IN1(n3264), .IN2(n3595), .IN3(elem08[14]), .IN4(n3262), .Q(
        n2858) );
  AO22X1 U1979 ( .IN1(n3264), .IN2(n3598), .IN3(elem08[15]), .IN4(n3262), .Q(
        n2859) );
  AO22X1 U1980 ( .IN1(n3264), .IN2(n3601), .IN3(elem08[16]), .IN4(n3262), .Q(
        n2860) );
  AO22X1 U1981 ( .IN1(n3264), .IN2(n3604), .IN3(elem08[17]), .IN4(n3262), .Q(
        n2861) );
  AO22X1 U1982 ( .IN1(n3264), .IN2(n3607), .IN3(elem08[18]), .IN4(n3262), .Q(
        n2862) );
  AO22X1 U1983 ( .IN1(n3265), .IN2(n3610), .IN3(elem08[19]), .IN4(n3262), .Q(
        n2863) );
  AO22X1 U1984 ( .IN1(n3264), .IN2(n3613), .IN3(elem08[20]), .IN4(n3261), .Q(
        n2864) );
  AO22X1 U1985 ( .IN1(n3265), .IN2(n3616), .IN3(elem08[21]), .IN4(n3261), .Q(
        n2865) );
  AO22X1 U1986 ( .IN1(n3264), .IN2(n3619), .IN3(elem08[22]), .IN4(n3261), .Q(
        n2866) );
  AO22X1 U1987 ( .IN1(n3265), .IN2(n3622), .IN3(elem08[23]), .IN4(n3261), .Q(
        n2867) );
  AO22X1 U1988 ( .IN1(n3264), .IN2(n3625), .IN3(elem08[24]), .IN4(n3261), .Q(
        n2868) );
  AO22X1 U1989 ( .IN1(n3265), .IN2(n3628), .IN3(elem08[25]), .IN4(n3261), .Q(
        n2869) );
  AO22X1 U1990 ( .IN1(n3265), .IN2(n3631), .IN3(elem08[26]), .IN4(n3261), .Q(
        n2870) );
  AO22X1 U1991 ( .IN1(n3265), .IN2(n3634), .IN3(elem08[27]), .IN4(n3261), .Q(
        n2871) );
  AO22X1 U1992 ( .IN1(n3265), .IN2(n3637), .IN3(elem08[28]), .IN4(n3261), .Q(
        n2872) );
  AO22X1 U1993 ( .IN1(n3265), .IN2(n3640), .IN3(elem08[29]), .IN4(n3261), .Q(
        n2873) );
  AO22X1 U1994 ( .IN1(n3265), .IN2(n3643), .IN3(elem08[30]), .IN4(n3261), .Q(
        n2874) );
  AO22X1 U1995 ( .IN1(n3265), .IN2(n3646), .IN3(elem08[31]), .IN4(n3261), .Q(
        n2875) );
  AND2X1 U1996 ( .IN1(n2248), .IN2(n2229), .Q(n2251) );
  AO22X1 U1997 ( .IN1(n2000), .IN2(n3552), .IN3(elem07[0]), .IN4(n2255), .Q(
        n2876) );
  AO22X1 U1998 ( .IN1(n2000), .IN2(n3555), .IN3(elem07[1]), .IN4(n2255), .Q(
        n2877) );
  AO22X1 U1999 ( .IN1(n2000), .IN2(n3558), .IN3(elem07[2]), .IN4(n2255), .Q(
        n2878) );
  AO22X1 U2000 ( .IN1(n2000), .IN2(n3561), .IN3(elem07[3]), .IN4(n2255), .Q(
        n2879) );
  AO22X1 U2001 ( .IN1(n2001), .IN2(n3564), .IN3(elem07[4]), .IN4(n2255), .Q(
        n2880) );
  AO22X1 U2002 ( .IN1(n3260), .IN2(n3567), .IN3(elem07[5]), .IN4(n2255), .Q(
        n2881) );
  AO22X1 U2003 ( .IN1(n3260), .IN2(n3570), .IN3(elem07[6]), .IN4(n2255), .Q(
        n2882) );
  AO22X1 U2004 ( .IN1(n2001), .IN2(n3573), .IN3(elem07[7]), .IN4(n2255), .Q(
        n2883) );
  AO22X1 U2005 ( .IN1(n3260), .IN2(n3576), .IN3(elem07[8]), .IN4(n1038), .Q(
        n2884) );
  AO22X1 U2006 ( .IN1(n3260), .IN2(n3579), .IN3(elem07[9]), .IN4(n1038), .Q(
        n2885) );
  AO22X1 U2007 ( .IN1(n2001), .IN2(n3582), .IN3(elem07[10]), .IN4(n1038), .Q(
        n2886) );
  AO22X1 U2008 ( .IN1(n2001), .IN2(n3585), .IN3(elem07[11]), .IN4(n1038), .Q(
        n2887) );
  AO22X1 U2009 ( .IN1(n2001), .IN2(n3589), .IN3(elem07[12]), .IN4(n1038), .Q(
        n2888) );
  AO22X1 U2010 ( .IN1(n2001), .IN2(n3592), .IN3(elem07[13]), .IN4(n1038), .Q(
        n2889) );
  AO22X1 U2011 ( .IN1(n2001), .IN2(n3595), .IN3(elem07[14]), .IN4(n1038), .Q(
        n2890) );
  AO22X1 U2012 ( .IN1(n2001), .IN2(n3598), .IN3(elem07[15]), .IN4(n1038), .Q(
        n2891) );
  AO22X1 U2013 ( .IN1(n2001), .IN2(n3601), .IN3(elem07[16]), .IN4(n1038), .Q(
        n2892) );
  AO22X1 U2014 ( .IN1(n2001), .IN2(n3604), .IN3(elem07[17]), .IN4(n1038), .Q(
        n2893) );
  AO22X1 U2015 ( .IN1(n2001), .IN2(n3607), .IN3(elem07[18]), .IN4(n1038), .Q(
        n2894) );
  AO22X1 U2016 ( .IN1(n3260), .IN2(n3610), .IN3(elem07[19]), .IN4(n1038), .Q(
        n2895) );
  AO22X1 U2017 ( .IN1(n2001), .IN2(n3613), .IN3(elem07[20]), .IN4(n1037), .Q(
        n2896) );
  AO22X1 U2018 ( .IN1(n3260), .IN2(n3616), .IN3(elem07[21]), .IN4(n1037), .Q(
        n2897) );
  AO22X1 U2019 ( .IN1(n2001), .IN2(n3619), .IN3(elem07[22]), .IN4(n1037), .Q(
        n2898) );
  AO22X1 U2020 ( .IN1(n3260), .IN2(n3622), .IN3(elem07[23]), .IN4(n1037), .Q(
        n2899) );
  AO22X1 U2021 ( .IN1(n2001), .IN2(n3625), .IN3(elem07[24]), .IN4(n1037), .Q(
        n2900) );
  AO22X1 U2022 ( .IN1(n3260), .IN2(n3628), .IN3(elem07[25]), .IN4(n1037), .Q(
        n2901) );
  AO22X1 U2023 ( .IN1(n3260), .IN2(n3631), .IN3(elem07[26]), .IN4(n1037), .Q(
        n2902) );
  AO22X1 U2024 ( .IN1(n3260), .IN2(n3634), .IN3(elem07[27]), .IN4(n1037), .Q(
        n2903) );
  AO22X1 U2025 ( .IN1(n3260), .IN2(n3637), .IN3(elem07[28]), .IN4(n1037), .Q(
        n2904) );
  AO22X1 U2026 ( .IN1(n3260), .IN2(n3640), .IN3(elem07[29]), .IN4(n1037), .Q(
        n2905) );
  AO22X1 U2027 ( .IN1(n3260), .IN2(n3643), .IN3(elem07[30]), .IN4(n1037), .Q(
        n2906) );
  AO22X1 U2028 ( .IN1(n3260), .IN2(n3646), .IN3(elem07[31]), .IN4(n1037), .Q(
        n2907) );
  AO22X1 U2029 ( .IN1(n1034), .IN2(n3552), .IN3(elem06[0]), .IN4(n2257), .Q(
        n2908) );
  AO22X1 U2030 ( .IN1(n1034), .IN2(n3555), .IN3(elem06[1]), .IN4(n2257), .Q(
        n2909) );
  AO22X1 U2031 ( .IN1(n1034), .IN2(n3558), .IN3(elem06[2]), .IN4(n2257), .Q(
        n2910) );
  AO22X1 U2032 ( .IN1(n1034), .IN2(n3561), .IN3(elem06[3]), .IN4(n2257), .Q(
        n2911) );
  AO22X1 U2033 ( .IN1(n1035), .IN2(n3564), .IN3(elem06[4]), .IN4(n2257), .Q(
        n2912) );
  AO22X1 U2034 ( .IN1(n1036), .IN2(n3567), .IN3(elem06[5]), .IN4(n2257), .Q(
        n2913) );
  AO22X1 U2035 ( .IN1(n1036), .IN2(n3570), .IN3(elem06[6]), .IN4(n2257), .Q(
        n2914) );
  AO22X1 U2036 ( .IN1(n1035), .IN2(n3573), .IN3(elem06[7]), .IN4(n2257), .Q(
        n2915) );
  AO22X1 U2037 ( .IN1(n1036), .IN2(n3576), .IN3(elem06[8]), .IN4(n1033), .Q(
        n2916) );
  AO22X1 U2038 ( .IN1(n1036), .IN2(n3579), .IN3(elem06[9]), .IN4(n1033), .Q(
        n2917) );
  AO22X1 U2039 ( .IN1(n1035), .IN2(n3582), .IN3(elem06[10]), .IN4(n1033), .Q(
        n2918) );
  AO22X1 U2040 ( .IN1(n1035), .IN2(n3585), .IN3(elem06[11]), .IN4(n1033), .Q(
        n2919) );
  AO22X1 U2041 ( .IN1(n1035), .IN2(n3589), .IN3(elem06[12]), .IN4(n1033), .Q(
        n2920) );
  AO22X1 U2042 ( .IN1(n1035), .IN2(n3592), .IN3(elem06[13]), .IN4(n1033), .Q(
        n2921) );
  AO22X1 U2043 ( .IN1(n1035), .IN2(n3595), .IN3(elem06[14]), .IN4(n1033), .Q(
        n2922) );
  AO22X1 U2044 ( .IN1(n1035), .IN2(n3598), .IN3(elem06[15]), .IN4(n1033), .Q(
        n2923) );
  AO22X1 U2045 ( .IN1(n1035), .IN2(n3601), .IN3(elem06[16]), .IN4(n1033), .Q(
        n2924) );
  AO22X1 U2046 ( .IN1(n1035), .IN2(n3604), .IN3(elem06[17]), .IN4(n1033), .Q(
        n2925) );
  AO22X1 U2047 ( .IN1(n1035), .IN2(n3607), .IN3(elem06[18]), .IN4(n1033), .Q(
        n2926) );
  AO22X1 U2048 ( .IN1(n1036), .IN2(n3610), .IN3(elem06[19]), .IN4(n1033), .Q(
        n2927) );
  AO22X1 U2049 ( .IN1(n1035), .IN2(n3613), .IN3(elem06[20]), .IN4(n1032), .Q(
        n2928) );
  AO22X1 U2050 ( .IN1(n1036), .IN2(n3616), .IN3(elem06[21]), .IN4(n1032), .Q(
        n2929) );
  AO22X1 U2051 ( .IN1(n1035), .IN2(n3619), .IN3(elem06[22]), .IN4(n1032), .Q(
        n2930) );
  AO22X1 U2052 ( .IN1(n1036), .IN2(n3622), .IN3(elem06[23]), .IN4(n1032), .Q(
        n2931) );
  AO22X1 U2053 ( .IN1(n1035), .IN2(n3625), .IN3(elem06[24]), .IN4(n1032), .Q(
        n2932) );
  AO22X1 U2054 ( .IN1(n1036), .IN2(n3628), .IN3(elem06[25]), .IN4(n1032), .Q(
        n2933) );
  AO22X1 U2055 ( .IN1(n1036), .IN2(n3631), .IN3(elem06[26]), .IN4(n1032), .Q(
        n2934) );
  AO22X1 U2056 ( .IN1(n1036), .IN2(n3634), .IN3(elem06[27]), .IN4(n1032), .Q(
        n2935) );
  AO22X1 U2057 ( .IN1(n1036), .IN2(n3637), .IN3(elem06[28]), .IN4(n1032), .Q(
        n2936) );
  AO22X1 U2058 ( .IN1(n1036), .IN2(n3640), .IN3(elem06[29]), .IN4(n1032), .Q(
        n2937) );
  AO22X1 U2059 ( .IN1(n1036), .IN2(n3643), .IN3(elem06[30]), .IN4(n1032), .Q(
        n2938) );
  AO22X1 U2060 ( .IN1(n1036), .IN2(n3646), .IN3(elem06[31]), .IN4(n1032), .Q(
        n2939) );
  AO22X1 U2061 ( .IN1(n1029), .IN2(n3552), .IN3(elem05[0]), .IN4(n2258), .Q(
        n2940) );
  AO22X1 U2062 ( .IN1(n1029), .IN2(n3555), .IN3(elem05[1]), .IN4(n2258), .Q(
        n2941) );
  AO22X1 U2063 ( .IN1(n1029), .IN2(n3558), .IN3(elem05[2]), .IN4(n2258), .Q(
        n2942) );
  AO22X1 U2064 ( .IN1(n1029), .IN2(n3561), .IN3(elem05[3]), .IN4(n2258), .Q(
        n2943) );
  AO22X1 U2065 ( .IN1(n1030), .IN2(n3564), .IN3(elem05[4]), .IN4(n2258), .Q(
        n2944) );
  AO22X1 U2066 ( .IN1(n1031), .IN2(n3567), .IN3(elem05[5]), .IN4(n2258), .Q(
        n2945) );
  AO22X1 U2067 ( .IN1(n1031), .IN2(n3570), .IN3(elem05[6]), .IN4(n2258), .Q(
        n2946) );
  AO22X1 U2068 ( .IN1(n1030), .IN2(n3573), .IN3(elem05[7]), .IN4(n2258), .Q(
        n2947) );
  AO22X1 U2069 ( .IN1(n1031), .IN2(n3576), .IN3(elem05[8]), .IN4(n1028), .Q(
        n2948) );
  AO22X1 U2070 ( .IN1(n1031), .IN2(n3579), .IN3(elem05[9]), .IN4(n1028), .Q(
        n2949) );
  AO22X1 U2071 ( .IN1(n1030), .IN2(n3582), .IN3(elem05[10]), .IN4(n1028), .Q(
        n2950) );
  AO22X1 U2072 ( .IN1(n1030), .IN2(n3585), .IN3(elem05[11]), .IN4(n1028), .Q(
        n2951) );
  AO22X1 U2073 ( .IN1(n1030), .IN2(n3589), .IN3(elem05[12]), .IN4(n1028), .Q(
        n2952) );
  AO22X1 U2074 ( .IN1(n1030), .IN2(n3592), .IN3(elem05[13]), .IN4(n1028), .Q(
        n2953) );
  AO22X1 U2075 ( .IN1(n1030), .IN2(n3595), .IN3(elem05[14]), .IN4(n1028), .Q(
        n2954) );
  AO22X1 U2076 ( .IN1(n1030), .IN2(n3598), .IN3(elem05[15]), .IN4(n1028), .Q(
        n2955) );
  AO22X1 U2077 ( .IN1(n1030), .IN2(n3601), .IN3(elem05[16]), .IN4(n1028), .Q(
        n2956) );
  AO22X1 U2078 ( .IN1(n1030), .IN2(n3604), .IN3(elem05[17]), .IN4(n1028), .Q(
        n2957) );
  AO22X1 U2079 ( .IN1(n1030), .IN2(n3607), .IN3(elem05[18]), .IN4(n1028), .Q(
        n2958) );
  AO22X1 U2080 ( .IN1(n1031), .IN2(n3610), .IN3(elem05[19]), .IN4(n1028), .Q(
        n2959) );
  AO22X1 U2081 ( .IN1(n1030), .IN2(n3613), .IN3(elem05[20]), .IN4(n1027), .Q(
        n2960) );
  AO22X1 U2082 ( .IN1(n1031), .IN2(n3616), .IN3(elem05[21]), .IN4(n1027), .Q(
        n2961) );
  AO22X1 U2083 ( .IN1(n1030), .IN2(n3619), .IN3(elem05[22]), .IN4(n1027), .Q(
        n2962) );
  AO22X1 U2084 ( .IN1(n1031), .IN2(n3622), .IN3(elem05[23]), .IN4(n1027), .Q(
        n2963) );
  AO22X1 U2085 ( .IN1(n1030), .IN2(n3625), .IN3(elem05[24]), .IN4(n1027), .Q(
        n2964) );
  AO22X1 U2086 ( .IN1(n1031), .IN2(n3628), .IN3(elem05[25]), .IN4(n1027), .Q(
        n2965) );
  AO22X1 U2087 ( .IN1(n1031), .IN2(n3631), .IN3(elem05[26]), .IN4(n1027), .Q(
        n2966) );
  AO22X1 U2088 ( .IN1(n1031), .IN2(n3634), .IN3(elem05[27]), .IN4(n1027), .Q(
        n2967) );
  AO22X1 U2089 ( .IN1(n1031), .IN2(n3637), .IN3(elem05[28]), .IN4(n1027), .Q(
        n2968) );
  AO22X1 U2090 ( .IN1(n1031), .IN2(n3640), .IN3(elem05[29]), .IN4(n1027), .Q(
        n2969) );
  AO22X1 U2091 ( .IN1(n1031), .IN2(n3643), .IN3(elem05[30]), .IN4(n1027), .Q(
        n2970) );
  AO22X1 U2092 ( .IN1(n1031), .IN2(n3646), .IN3(elem05[31]), .IN4(n1027), .Q(
        n2971) );
  AO22X1 U2093 ( .IN1(n1024), .IN2(n3552), .IN3(elem04[0]), .IN4(n2259), .Q(
        n2972) );
  AO22X1 U2094 ( .IN1(n1024), .IN2(n3555), .IN3(elem04[1]), .IN4(n2259), .Q(
        n2973) );
  AO22X1 U2095 ( .IN1(n1024), .IN2(n3558), .IN3(elem04[2]), .IN4(n2259), .Q(
        n2974) );
  AO22X1 U2096 ( .IN1(n1024), .IN2(n3561), .IN3(elem04[3]), .IN4(n2259), .Q(
        n2975) );
  AO22X1 U2097 ( .IN1(n1025), .IN2(n3564), .IN3(elem04[4]), .IN4(n2259), .Q(
        n2976) );
  AO22X1 U2098 ( .IN1(n1026), .IN2(n3567), .IN3(elem04[5]), .IN4(n2259), .Q(
        n2977) );
  AO22X1 U2099 ( .IN1(n1026), .IN2(n3570), .IN3(elem04[6]), .IN4(n2259), .Q(
        n2978) );
  AO22X1 U2100 ( .IN1(n1025), .IN2(n3573), .IN3(elem04[7]), .IN4(n2259), .Q(
        n2979) );
  AO22X1 U2101 ( .IN1(n1026), .IN2(n3576), .IN3(elem04[8]), .IN4(n1023), .Q(
        n2980) );
  AO22X1 U2102 ( .IN1(n1026), .IN2(n3579), .IN3(elem04[9]), .IN4(n1023), .Q(
        n2981) );
  AO22X1 U2103 ( .IN1(n1025), .IN2(n3582), .IN3(elem04[10]), .IN4(n1023), .Q(
        n2982) );
  AO22X1 U2104 ( .IN1(n1025), .IN2(n3585), .IN3(elem04[11]), .IN4(n1023), .Q(
        n2983) );
  AO22X1 U2105 ( .IN1(n1025), .IN2(n3590), .IN3(elem04[12]), .IN4(n1023), .Q(
        n2984) );
  AO22X1 U2106 ( .IN1(n1025), .IN2(n3593), .IN3(elem04[13]), .IN4(n1023), .Q(
        n2985) );
  AO22X1 U2107 ( .IN1(n1025), .IN2(n3596), .IN3(elem04[14]), .IN4(n1023), .Q(
        n2986) );
  AO22X1 U2108 ( .IN1(n1025), .IN2(n3599), .IN3(elem04[15]), .IN4(n1023), .Q(
        n2987) );
  AO22X1 U2109 ( .IN1(n1025), .IN2(n3602), .IN3(elem04[16]), .IN4(n1023), .Q(
        n2988) );
  AO22X1 U2110 ( .IN1(n1025), .IN2(n3605), .IN3(elem04[17]), .IN4(n1023), .Q(
        n2989) );
  AO22X1 U2111 ( .IN1(n1025), .IN2(n3608), .IN3(elem04[18]), .IN4(n1023), .Q(
        n2990) );
  AO22X1 U2112 ( .IN1(n1026), .IN2(n3611), .IN3(elem04[19]), .IN4(n1023), .Q(
        n2991) );
  AO22X1 U2113 ( .IN1(n1025), .IN2(n3614), .IN3(elem04[20]), .IN4(n1022), .Q(
        n2992) );
  AO22X1 U2114 ( .IN1(n1026), .IN2(n3617), .IN3(elem04[21]), .IN4(n1022), .Q(
        n2993) );
  AO22X1 U2115 ( .IN1(n1025), .IN2(n3620), .IN3(elem04[22]), .IN4(n1022), .Q(
        n2994) );
  AO22X1 U2116 ( .IN1(n1026), .IN2(n3623), .IN3(elem04[23]), .IN4(n1022), .Q(
        n2995) );
  AO22X1 U2117 ( .IN1(n1025), .IN2(n3626), .IN3(elem04[24]), .IN4(n1022), .Q(
        n2996) );
  AO22X1 U2118 ( .IN1(n1026), .IN2(n3629), .IN3(elem04[25]), .IN4(n1022), .Q(
        n2997) );
  AO22X1 U2119 ( .IN1(n1026), .IN2(n3632), .IN3(elem04[26]), .IN4(n1022), .Q(
        n2998) );
  AO22X1 U2120 ( .IN1(n1026), .IN2(n3635), .IN3(elem04[27]), .IN4(n1022), .Q(
        n2999) );
  AO22X1 U2121 ( .IN1(n1026), .IN2(n3638), .IN3(elem04[28]), .IN4(n1022), .Q(
        n3000) );
  AO22X1 U2122 ( .IN1(n1026), .IN2(n3641), .IN3(elem04[29]), .IN4(n1022), .Q(
        n3001) );
  AO22X1 U2123 ( .IN1(n1026), .IN2(n3644), .IN3(elem04[30]), .IN4(n1022), .Q(
        n3002) );
  AO22X1 U2124 ( .IN1(n1026), .IN2(n3647), .IN3(elem04[31]), .IN4(n1022), .Q(
        n3003) );
  AND2X1 U2125 ( .IN1(n2248), .IN2(n2236), .Q(n2256) );
  AO22X1 U2126 ( .IN1(n1021), .IN2(n3553), .IN3(elem03[0]), .IN4(n2260), .Q(
        n3004) );
  AO22X1 U2127 ( .IN1(n1020), .IN2(n3556), .IN3(elem03[1]), .IN4(n2260), .Q(
        n3005) );
  AO22X1 U2128 ( .IN1(n1021), .IN2(n3559), .IN3(elem03[2]), .IN4(n2260), .Q(
        n3006) );
  AO22X1 U2129 ( .IN1(n1020), .IN2(n3562), .IN3(elem03[3]), .IN4(n2260), .Q(
        n3007) );
  AO22X1 U2130 ( .IN1(n1020), .IN2(n3565), .IN3(elem03[4]), .IN4(n2260), .Q(
        n3008) );
  AO22X1 U2131 ( .IN1(n1021), .IN2(n3568), .IN3(elem03[5]), .IN4(n2260), .Q(
        n3009) );
  AO22X1 U2132 ( .IN1(n1021), .IN2(n3571), .IN3(elem03[6]), .IN4(n2260), .Q(
        n3010) );
  AO22X1 U2133 ( .IN1(n1020), .IN2(n3574), .IN3(elem03[7]), .IN4(n2260), .Q(
        n3011) );
  AO22X1 U2134 ( .IN1(n1021), .IN2(n3577), .IN3(elem03[8]), .IN4(n1019), .Q(
        n3012) );
  AO22X1 U2135 ( .IN1(n1021), .IN2(n3580), .IN3(elem03[9]), .IN4(n1019), .Q(
        n3013) );
  AO22X1 U2136 ( .IN1(n1020), .IN2(n3583), .IN3(elem03[10]), .IN4(n1019), .Q(
        n3014) );
  AO22X1 U2137 ( .IN1(n1020), .IN2(n3586), .IN3(elem03[11]), .IN4(n1019), .Q(
        n3015) );
  AO22X1 U2138 ( .IN1(n1020), .IN2(n3590), .IN3(elem03[12]), .IN4(n1019), .Q(
        n3016) );
  AO22X1 U2139 ( .IN1(n1020), .IN2(n3593), .IN3(elem03[13]), .IN4(n1019), .Q(
        n3017) );
  AO22X1 U2140 ( .IN1(n1020), .IN2(n3596), .IN3(elem03[14]), .IN4(n1019), .Q(
        n3018) );
  AO22X1 U2141 ( .IN1(n1020), .IN2(n3599), .IN3(elem03[15]), .IN4(n1019), .Q(
        n3019) );
  AO22X1 U2142 ( .IN1(n1020), .IN2(n3602), .IN3(elem03[16]), .IN4(n1019), .Q(
        n3020) );
  AO22X1 U2143 ( .IN1(n1020), .IN2(n3605), .IN3(elem03[17]), .IN4(n1019), .Q(
        n3021) );
  AO22X1 U2144 ( .IN1(n1020), .IN2(n3608), .IN3(elem03[18]), .IN4(n1019), .Q(
        n3022) );
  AO22X1 U2145 ( .IN1(n1021), .IN2(n3611), .IN3(elem03[19]), .IN4(n1019), .Q(
        n3023) );
  AO22X1 U2146 ( .IN1(n1020), .IN2(n3614), .IN3(elem03[20]), .IN4(n1018), .Q(
        n3024) );
  AO22X1 U2147 ( .IN1(n1021), .IN2(n3617), .IN3(elem03[21]), .IN4(n1018), .Q(
        n3025) );
  AO22X1 U2148 ( .IN1(n1020), .IN2(n3620), .IN3(elem03[22]), .IN4(n1018), .Q(
        n3026) );
  AO22X1 U2149 ( .IN1(n1021), .IN2(n3623), .IN3(elem03[23]), .IN4(n1018), .Q(
        n3027) );
  AO22X1 U2150 ( .IN1(n1020), .IN2(n3626), .IN3(elem03[24]), .IN4(n1018), .Q(
        n3028) );
  AO22X1 U2151 ( .IN1(n1021), .IN2(n3629), .IN3(elem03[25]), .IN4(n1018), .Q(
        n3029) );
  AO22X1 U2152 ( .IN1(n1021), .IN2(n3632), .IN3(elem03[26]), .IN4(n1018), .Q(
        n3030) );
  AO22X1 U2153 ( .IN1(n1021), .IN2(n3635), .IN3(elem03[27]), .IN4(n1018), .Q(
        n3031) );
  AO22X1 U2154 ( .IN1(n1021), .IN2(n3638), .IN3(elem03[28]), .IN4(n1018), .Q(
        n3032) );
  AO22X1 U2155 ( .IN1(n1021), .IN2(n3641), .IN3(elem03[29]), .IN4(n1018), .Q(
        n3033) );
  AO22X1 U2156 ( .IN1(n1021), .IN2(n3644), .IN3(elem03[30]), .IN4(n1018), .Q(
        n3034) );
  AO22X1 U2157 ( .IN1(n1021), .IN2(n3647), .IN3(elem03[31]), .IN4(n1018), .Q(
        n3035) );
  AO22X1 U2158 ( .IN1(n1017), .IN2(n3552), .IN3(elem02[0]), .IN4(n2262), .Q(
        n3036) );
  AO22X1 U2159 ( .IN1(n1016), .IN2(n3555), .IN3(elem02[1]), .IN4(n2262), .Q(
        n3037) );
  AO22X1 U2160 ( .IN1(n1017), .IN2(n3558), .IN3(elem02[2]), .IN4(n2262), .Q(
        n3038) );
  AO22X1 U2161 ( .IN1(n1016), .IN2(n3561), .IN3(elem02[3]), .IN4(n2262), .Q(
        n3039) );
  AO22X1 U2162 ( .IN1(n1016), .IN2(n3564), .IN3(elem02[4]), .IN4(n2262), .Q(
        n3040) );
  AO22X1 U2163 ( .IN1(n1017), .IN2(n3567), .IN3(elem02[5]), .IN4(n2262), .Q(
        n3041) );
  AO22X1 U2164 ( .IN1(n1017), .IN2(n3570), .IN3(elem02[6]), .IN4(n2262), .Q(
        n3042) );
  AO22X1 U2165 ( .IN1(n1016), .IN2(n3573), .IN3(elem02[7]), .IN4(n2262), .Q(
        n3043) );
  AO22X1 U2166 ( .IN1(n1017), .IN2(n3576), .IN3(elem02[8]), .IN4(n1015), .Q(
        n3044) );
  AO22X1 U2167 ( .IN1(n1017), .IN2(n3579), .IN3(elem02[9]), .IN4(n1015), .Q(
        n3045) );
  AO22X1 U2168 ( .IN1(n1016), .IN2(n3582), .IN3(elem02[10]), .IN4(n1015), .Q(
        n3046) );
  AO22X1 U2169 ( .IN1(n1016), .IN2(n3585), .IN3(elem02[11]), .IN4(n1015), .Q(
        n3047) );
  AO22X1 U2170 ( .IN1(n1016), .IN2(n3590), .IN3(elem02[12]), .IN4(n1015), .Q(
        n3048) );
  AO22X1 U2171 ( .IN1(n1016), .IN2(n3593), .IN3(elem02[13]), .IN4(n1015), .Q(
        n3049) );
  AO22X1 U2172 ( .IN1(n1016), .IN2(n3596), .IN3(elem02[14]), .IN4(n1015), .Q(
        n3050) );
  AO22X1 U2173 ( .IN1(n1016), .IN2(n3599), .IN3(elem02[15]), .IN4(n1015), .Q(
        n3051) );
  AO22X1 U2174 ( .IN1(n1016), .IN2(n3602), .IN3(elem02[16]), .IN4(n1015), .Q(
        n3052) );
  AO22X1 U2175 ( .IN1(n1016), .IN2(n3605), .IN3(elem02[17]), .IN4(n1015), .Q(
        n3053) );
  AO22X1 U2176 ( .IN1(n1016), .IN2(n3608), .IN3(elem02[18]), .IN4(n1015), .Q(
        n3054) );
  AO22X1 U2177 ( .IN1(n1017), .IN2(n3611), .IN3(elem02[19]), .IN4(n1015), .Q(
        n3055) );
  AO22X1 U2178 ( .IN1(n1016), .IN2(n3614), .IN3(elem02[20]), .IN4(n1014), .Q(
        n3056) );
  AO22X1 U2179 ( .IN1(n1017), .IN2(n3617), .IN3(elem02[21]), .IN4(n1014), .Q(
        n3057) );
  AO22X1 U2180 ( .IN1(n1016), .IN2(n3620), .IN3(elem02[22]), .IN4(n1014), .Q(
        n3058) );
  AO22X1 U2181 ( .IN1(n1017), .IN2(n3623), .IN3(elem02[23]), .IN4(n1014), .Q(
        n3059) );
  AO22X1 U2182 ( .IN1(n1016), .IN2(n3626), .IN3(elem02[24]), .IN4(n1014), .Q(
        n3060) );
  AO22X1 U2183 ( .IN1(n1017), .IN2(n3629), .IN3(elem02[25]), .IN4(n1014), .Q(
        n3061) );
  AO22X1 U2184 ( .IN1(n1017), .IN2(n3632), .IN3(elem02[26]), .IN4(n1014), .Q(
        n3062) );
  AO22X1 U2185 ( .IN1(n1017), .IN2(n3635), .IN3(elem02[27]), .IN4(n1014), .Q(
        n3063) );
  AO22X1 U2186 ( .IN1(n1017), .IN2(n3638), .IN3(elem02[28]), .IN4(n1014), .Q(
        n3064) );
  AO22X1 U2187 ( .IN1(n1017), .IN2(n3641), .IN3(elem02[29]), .IN4(n1014), .Q(
        n3065) );
  AO22X1 U2188 ( .IN1(n1017), .IN2(n3644), .IN3(elem02[30]), .IN4(n1014), .Q(
        n3066) );
  AO22X1 U2189 ( .IN1(n1017), .IN2(n3647), .IN3(elem02[31]), .IN4(n1014), .Q(
        n3067) );
  AO22X1 U2190 ( .IN1(n1013), .IN2(n3552), .IN3(elem01[0]), .IN4(n2263), .Q(
        n3068) );
  AO22X1 U2191 ( .IN1(n1012), .IN2(n3555), .IN3(elem01[1]), .IN4(n2263), .Q(
        n3069) );
  AO22X1 U2192 ( .IN1(n1013), .IN2(n3558), .IN3(elem01[2]), .IN4(n2263), .Q(
        n3070) );
  AO22X1 U2193 ( .IN1(n1012), .IN2(n3561), .IN3(elem01[3]), .IN4(n2263), .Q(
        n3071) );
  AO22X1 U2194 ( .IN1(n1012), .IN2(n3564), .IN3(elem01[4]), .IN4(n2263), .Q(
        n3072) );
  AO22X1 U2195 ( .IN1(n1013), .IN2(n3567), .IN3(elem01[5]), .IN4(n2263), .Q(
        n3073) );
  AO22X1 U2196 ( .IN1(n1013), .IN2(n3570), .IN3(elem01[6]), .IN4(n2263), .Q(
        n3074) );
  AO22X1 U2197 ( .IN1(n1012), .IN2(n3573), .IN3(elem01[7]), .IN4(n2263), .Q(
        n3075) );
  AO22X1 U2198 ( .IN1(n1013), .IN2(n3576), .IN3(elem01[8]), .IN4(n1011), .Q(
        n3076) );
  AO22X1 U2199 ( .IN1(n1013), .IN2(n3579), .IN3(elem01[9]), .IN4(n1011), .Q(
        n3077) );
  AO22X1 U2200 ( .IN1(n1012), .IN2(n3582), .IN3(elem01[10]), .IN4(n1011), .Q(
        n3078) );
  AO22X1 U2201 ( .IN1(n1012), .IN2(n3585), .IN3(elem01[11]), .IN4(n1011), .Q(
        n3079) );
  AO22X1 U2202 ( .IN1(n1012), .IN2(n3590), .IN3(elem01[12]), .IN4(n1011), .Q(
        n3080) );
  AO22X1 U2203 ( .IN1(n1012), .IN2(n3593), .IN3(elem01[13]), .IN4(n1011), .Q(
        n3081) );
  AO22X1 U2204 ( .IN1(n1012), .IN2(n3596), .IN3(elem01[14]), .IN4(n1011), .Q(
        n3082) );
  AO22X1 U2205 ( .IN1(n1012), .IN2(n3599), .IN3(elem01[15]), .IN4(n1011), .Q(
        n3083) );
  AO22X1 U2206 ( .IN1(n1012), .IN2(n3602), .IN3(elem01[16]), .IN4(n1011), .Q(
        n3084) );
  AO22X1 U2207 ( .IN1(n1012), .IN2(n3605), .IN3(elem01[17]), .IN4(n1011), .Q(
        n3085) );
  AO22X1 U2208 ( .IN1(n1012), .IN2(n3608), .IN3(elem01[18]), .IN4(n1011), .Q(
        n3086) );
  AO22X1 U2209 ( .IN1(n1013), .IN2(n3611), .IN3(elem01[19]), .IN4(n1011), .Q(
        n3087) );
  AO22X1 U2210 ( .IN1(n1012), .IN2(n3614), .IN3(elem01[20]), .IN4(n1010), .Q(
        n3088) );
  AO22X1 U2211 ( .IN1(n1013), .IN2(n3617), .IN3(elem01[21]), .IN4(n1010), .Q(
        n3089) );
  AO22X1 U2212 ( .IN1(n1012), .IN2(n3620), .IN3(elem01[22]), .IN4(n1010), .Q(
        n3090) );
  AO22X1 U2213 ( .IN1(n1013), .IN2(n3623), .IN3(elem01[23]), .IN4(n1010), .Q(
        n3091) );
  AO22X1 U2214 ( .IN1(n1012), .IN2(n3626), .IN3(elem01[24]), .IN4(n1010), .Q(
        n3092) );
  AO22X1 U2215 ( .IN1(n1013), .IN2(n3629), .IN3(elem01[25]), .IN4(n1010), .Q(
        n3093) );
  AO22X1 U2216 ( .IN1(n1013), .IN2(n3632), .IN3(elem01[26]), .IN4(n1010), .Q(
        n3094) );
  AO22X1 U2217 ( .IN1(n1013), .IN2(n3635), .IN3(elem01[27]), .IN4(n1010), .Q(
        n3095) );
  AO22X1 U2218 ( .IN1(n1013), .IN2(n3638), .IN3(elem01[28]), .IN4(n1010), .Q(
        n3096) );
  AO22X1 U2219 ( .IN1(n1013), .IN2(n3641), .IN3(elem01[29]), .IN4(n1010), .Q(
        n3097) );
  AO22X1 U2220 ( .IN1(n1013), .IN2(n3644), .IN3(elem01[30]), .IN4(n1010), .Q(
        n3098) );
  AO22X1 U2221 ( .IN1(n1013), .IN2(n3647), .IN3(elem01[31]), .IN4(n1010), .Q(
        n3099) );
  AND2X1 U2222 ( .IN1(n2248), .IN2(n2242), .Q(n2261) );
  AO22X1 U2223 ( .IN1(n1008), .IN2(n3552), .IN3(elem31[0]), .IN4(n2264), .Q(
        n3100) );
  AO22X1 U2224 ( .IN1(n1007), .IN2(n3555), .IN3(elem31[1]), .IN4(n1006), .Q(
        n3101) );
  AO22X1 U2225 ( .IN1(n1007), .IN2(n3558), .IN3(elem31[2]), .IN4(n2264), .Q(
        n3102) );
  AO22X1 U2226 ( .IN1(n1007), .IN2(n3561), .IN3(elem31[3]), .IN4(n2264), .Q(
        n3103) );
  AO22X1 U2227 ( .IN1(n1007), .IN2(n3564), .IN3(elem31[4]), .IN4(n2264), .Q(
        n3104) );
  AO22X1 U2228 ( .IN1(n1009), .IN2(n3567), .IN3(elem31[5]), .IN4(n2264), .Q(
        n3105) );
  AO22X1 U2229 ( .IN1(n1008), .IN2(n3570), .IN3(elem31[6]), .IN4(n2264), .Q(
        n3106) );
  AO22X1 U2230 ( .IN1(n1007), .IN2(n3573), .IN3(elem31[7]), .IN4(n2264), .Q(
        n3107) );
  AO22X1 U2231 ( .IN1(n1009), .IN2(n3576), .IN3(elem31[8]), .IN4(n1006), .Q(
        n3108) );
  AO22X1 U2232 ( .IN1(n1008), .IN2(n3579), .IN3(elem31[9]), .IN4(n1006), .Q(
        n3109) );
  AO22X1 U2233 ( .IN1(n1007), .IN2(n3582), .IN3(elem31[10]), .IN4(n1006), .Q(
        n3110) );
  AO22X1 U2234 ( .IN1(n1007), .IN2(n3585), .IN3(elem31[11]), .IN4(n1006), .Q(
        n3111) );
  AO22X1 U2235 ( .IN1(n1007), .IN2(n3590), .IN3(elem31[12]), .IN4(n1006), .Q(
        n3112) );
  AO22X1 U2236 ( .IN1(n1007), .IN2(n3593), .IN3(elem31[13]), .IN4(n1006), .Q(
        n3113) );
  AO22X1 U2237 ( .IN1(n1007), .IN2(n3596), .IN3(elem31[14]), .IN4(n1006), .Q(
        n3114) );
  AO22X1 U2238 ( .IN1(n1007), .IN2(n3599), .IN3(elem31[15]), .IN4(n1006), .Q(
        n3115) );
  AO22X1 U2239 ( .IN1(n1007), .IN2(n3602), .IN3(elem31[16]), .IN4(n1006), .Q(
        n3116) );
  AO22X1 U2240 ( .IN1(n1007), .IN2(n3605), .IN3(elem31[17]), .IN4(n1006), .Q(
        n3117) );
  AO22X1 U2241 ( .IN1(n1008), .IN2(n3608), .IN3(elem31[18]), .IN4(n1006), .Q(
        n3118) );
  AO22X1 U2242 ( .IN1(n1008), .IN2(n3611), .IN3(elem31[19]), .IN4(n1006), .Q(
        n3119) );
  AO22X1 U2243 ( .IN1(n1008), .IN2(n3614), .IN3(elem31[20]), .IN4(n1005), .Q(
        n3120) );
  AO22X1 U2244 ( .IN1(n1008), .IN2(n3617), .IN3(elem31[21]), .IN4(n1005), .Q(
        n3121) );
  AO22X1 U2245 ( .IN1(n1008), .IN2(n3620), .IN3(elem31[22]), .IN4(n1005), .Q(
        n3122) );
  AO22X1 U2246 ( .IN1(n1008), .IN2(n3623), .IN3(elem31[23]), .IN4(n1005), .Q(
        n3123) );
  AO22X1 U2247 ( .IN1(n1008), .IN2(n3626), .IN3(elem31[24]), .IN4(n1005), .Q(
        n3124) );
  AO22X1 U2248 ( .IN1(n1009), .IN2(n3629), .IN3(elem31[25]), .IN4(n1005), .Q(
        n3125) );
  AO22X1 U2249 ( .IN1(n1009), .IN2(n3632), .IN3(elem31[26]), .IN4(n1005), .Q(
        n3126) );
  AO22X1 U2250 ( .IN1(n1009), .IN2(n3635), .IN3(elem31[27]), .IN4(n1005), .Q(
        n3127) );
  AO22X1 U2251 ( .IN1(n1009), .IN2(n3638), .IN3(elem31[28]), .IN4(n1005), .Q(
        n3128) );
  AO22X1 U2252 ( .IN1(n1009), .IN2(n3641), .IN3(elem31[29]), .IN4(n1005), .Q(
        n3129) );
  AO22X1 U2253 ( .IN1(n1009), .IN2(n3644), .IN3(elem31[30]), .IN4(n1005), .Q(
        n3130) );
  AO22X1 U2254 ( .IN1(n1009), .IN2(n3647), .IN3(elem31[31]), .IN4(n1005), .Q(
        n3131) );
  AO22X1 U2255 ( .IN1(n1002), .IN2(n3552), .IN3(elem28[0]), .IN4(n2266), .Q(
        n3132) );
  AO22X1 U2256 ( .IN1(n1002), .IN2(n3555), .IN3(elem28[1]), .IN4(n2266), .Q(
        n3133) );
  AO22X1 U2257 ( .IN1(n1002), .IN2(n3558), .IN3(elem28[2]), .IN4(n2266), .Q(
        n3134) );
  AO22X1 U2258 ( .IN1(n1002), .IN2(n3561), .IN3(elem28[3]), .IN4(n2266), .Q(
        n3135) );
  AO22X1 U2259 ( .IN1(n1003), .IN2(n3564), .IN3(elem28[4]), .IN4(n2266), .Q(
        n3136) );
  AO22X1 U2260 ( .IN1(n1004), .IN2(n3567), .IN3(elem28[5]), .IN4(n2266), .Q(
        n3137) );
  AO22X1 U2261 ( .IN1(n1004), .IN2(n3570), .IN3(elem28[6]), .IN4(n2266), .Q(
        n3138) );
  AO22X1 U2262 ( .IN1(n1003), .IN2(n3573), .IN3(elem28[7]), .IN4(n2266), .Q(
        n3139) );
  AO22X1 U2263 ( .IN1(n1004), .IN2(n3576), .IN3(elem28[8]), .IN4(n1001), .Q(
        n3140) );
  AO22X1 U2264 ( .IN1(n1004), .IN2(n3579), .IN3(elem28[9]), .IN4(n1001), .Q(
        n3141) );
  AO22X1 U2265 ( .IN1(n1003), .IN2(n3582), .IN3(elem28[10]), .IN4(n1001), .Q(
        n3142) );
  AO22X1 U2266 ( .IN1(n1003), .IN2(n3585), .IN3(elem28[11]), .IN4(n1001), .Q(
        n3143) );
  AO22X1 U2267 ( .IN1(n1003), .IN2(n3590), .IN3(elem28[12]), .IN4(n1001), .Q(
        n3144) );
  AO22X1 U2268 ( .IN1(n1003), .IN2(n3593), .IN3(elem28[13]), .IN4(n1001), .Q(
        n3145) );
  AO22X1 U2269 ( .IN1(n1003), .IN2(n3596), .IN3(elem28[14]), .IN4(n1001), .Q(
        n3146) );
  AO22X1 U2270 ( .IN1(n1003), .IN2(n3599), .IN3(elem28[15]), .IN4(n1001), .Q(
        n3147) );
  AO22X1 U2271 ( .IN1(n1003), .IN2(n3602), .IN3(elem28[16]), .IN4(n1001), .Q(
        n3148) );
  AO22X1 U2272 ( .IN1(n1003), .IN2(n3605), .IN3(elem28[17]), .IN4(n1001), .Q(
        n3149) );
  AO22X1 U2273 ( .IN1(n1003), .IN2(n3608), .IN3(elem28[18]), .IN4(n1001), .Q(
        n3150) );
  AO22X1 U2274 ( .IN1(n1004), .IN2(n3611), .IN3(elem28[19]), .IN4(n1001), .Q(
        n3151) );
  AO22X1 U2275 ( .IN1(n1003), .IN2(n3614), .IN3(elem28[20]), .IN4(n1000), .Q(
        n3152) );
  AO22X1 U2276 ( .IN1(n1004), .IN2(n3617), .IN3(elem28[21]), .IN4(n1000), .Q(
        n3153) );
  AO22X1 U2277 ( .IN1(n1003), .IN2(n3620), .IN3(elem28[22]), .IN4(n1000), .Q(
        n3154) );
  AO22X1 U2278 ( .IN1(n1004), .IN2(n3623), .IN3(elem28[23]), .IN4(n1000), .Q(
        n3155) );
  AO22X1 U2279 ( .IN1(n1003), .IN2(n3626), .IN3(elem28[24]), .IN4(n1000), .Q(
        n3156) );
  AO22X1 U2280 ( .IN1(n1004), .IN2(n3629), .IN3(elem28[25]), .IN4(n1000), .Q(
        n3157) );
  AO22X1 U2281 ( .IN1(n1004), .IN2(n3632), .IN3(elem28[26]), .IN4(n1000), .Q(
        n3158) );
  AO22X1 U2282 ( .IN1(n1004), .IN2(n3635), .IN3(elem28[27]), .IN4(n1000), .Q(
        n3159) );
  AO22X1 U2283 ( .IN1(n1004), .IN2(n3638), .IN3(elem28[28]), .IN4(n1000), .Q(
        n3160) );
  AO22X1 U2284 ( .IN1(n1004), .IN2(n3641), .IN3(elem28[29]), .IN4(n1000), .Q(
        n3161) );
  AO22X1 U2285 ( .IN1(n1004), .IN2(n3644), .IN3(elem28[30]), .IN4(n1000), .Q(
        n3162) );
  AO22X1 U2286 ( .IN1(n1004), .IN2(n3647), .IN3(elem28[31]), .IN4(n1000), .Q(
        n3163) );
  AO22X1 U2287 ( .IN1(n998), .IN2(n3552), .IN3(elem29[0]), .IN4(n2267), .Q(
        n3164) );
  AO22X1 U2288 ( .IN1(n997), .IN2(n3555), .IN3(elem29[1]), .IN4(n996), .Q(
        n3165) );
  AO22X1 U2289 ( .IN1(n997), .IN2(n3558), .IN3(elem29[2]), .IN4(n2267), .Q(
        n3166) );
  AO22X1 U2290 ( .IN1(n997), .IN2(n3561), .IN3(elem29[3]), .IN4(n2267), .Q(
        n3167) );
  AO22X1 U2291 ( .IN1(n997), .IN2(n3564), .IN3(elem29[4]), .IN4(n2267), .Q(
        n3168) );
  AO22X1 U2292 ( .IN1(n999), .IN2(n3567), .IN3(elem29[5]), .IN4(n2267), .Q(
        n3169) );
  AO22X1 U2293 ( .IN1(n998), .IN2(n3570), .IN3(elem29[6]), .IN4(n2267), .Q(
        n3170) );
  AO22X1 U2294 ( .IN1(n997), .IN2(n3573), .IN3(elem29[7]), .IN4(n2267), .Q(
        n3171) );
  AO22X1 U2295 ( .IN1(n999), .IN2(n3576), .IN3(elem29[8]), .IN4(n996), .Q(
        n3172) );
  AO22X1 U2296 ( .IN1(n998), .IN2(n3579), .IN3(elem29[9]), .IN4(n996), .Q(
        n3173) );
  AO22X1 U2297 ( .IN1(n997), .IN2(n3582), .IN3(elem29[10]), .IN4(n996), .Q(
        n3174) );
  AO22X1 U2298 ( .IN1(n997), .IN2(n3585), .IN3(elem29[11]), .IN4(n996), .Q(
        n3175) );
  AO22X1 U2299 ( .IN1(n997), .IN2(n3590), .IN3(elem29[12]), .IN4(n996), .Q(
        n3176) );
  AO22X1 U2300 ( .IN1(n997), .IN2(n3593), .IN3(elem29[13]), .IN4(n996), .Q(
        n3177) );
  AO22X1 U2301 ( .IN1(n997), .IN2(n3596), .IN3(elem29[14]), .IN4(n996), .Q(
        n3178) );
  AO22X1 U2302 ( .IN1(n997), .IN2(n3599), .IN3(elem29[15]), .IN4(n996), .Q(
        n3179) );
  AO22X1 U2303 ( .IN1(n997), .IN2(n3602), .IN3(elem29[16]), .IN4(n996), .Q(
        n3180) );
  AO22X1 U2304 ( .IN1(n997), .IN2(n3605), .IN3(elem29[17]), .IN4(n996), .Q(
        n3181) );
  AO22X1 U2305 ( .IN1(n998), .IN2(n3608), .IN3(elem29[18]), .IN4(n996), .Q(
        n3182) );
  AO22X1 U2306 ( .IN1(n998), .IN2(n3611), .IN3(elem29[19]), .IN4(n996), .Q(
        n3183) );
  AO22X1 U2307 ( .IN1(n998), .IN2(n3614), .IN3(elem29[20]), .IN4(n995), .Q(
        n3184) );
  AO22X1 U2308 ( .IN1(n998), .IN2(n3617), .IN3(elem29[21]), .IN4(n995), .Q(
        n3185) );
  AO22X1 U2309 ( .IN1(n998), .IN2(n3620), .IN3(elem29[22]), .IN4(n995), .Q(
        n3186) );
  AO22X1 U2310 ( .IN1(n998), .IN2(n3623), .IN3(elem29[23]), .IN4(n995), .Q(
        n3187) );
  AO22X1 U2311 ( .IN1(n998), .IN2(n3626), .IN3(elem29[24]), .IN4(n995), .Q(
        n3188) );
  AO22X1 U2312 ( .IN1(n999), .IN2(n3629), .IN3(elem29[25]), .IN4(n995), .Q(
        n3189) );
  AO22X1 U2313 ( .IN1(n999), .IN2(n3632), .IN3(elem29[26]), .IN4(n995), .Q(
        n3190) );
  AO22X1 U2314 ( .IN1(n999), .IN2(n3635), .IN3(elem29[27]), .IN4(n995), .Q(
        n3191) );
  AO22X1 U2315 ( .IN1(n999), .IN2(n3638), .IN3(elem29[28]), .IN4(n995), .Q(
        n3192) );
  AO22X1 U2316 ( .IN1(n999), .IN2(n3641), .IN3(elem29[29]), .IN4(n995), .Q(
        n3193) );
  AO22X1 U2317 ( .IN1(n999), .IN2(n3644), .IN3(elem29[30]), .IN4(n995), .Q(
        n3194) );
  AO22X1 U2318 ( .IN1(n999), .IN2(n3647), .IN3(elem29[31]), .IN4(n995), .Q(
        n3195) );
  AO22X1 U2319 ( .IN1(n3552), .IN2(n3364), .IN3(elem30[0]), .IN4(n3361), .Q(
        n3196) );
  AO22X1 U2320 ( .IN1(n3555), .IN2(n3364), .IN3(elem30[1]), .IN4(n3361), .Q(
        n3197) );
  AO22X1 U2321 ( .IN1(n3558), .IN2(n3364), .IN3(elem30[2]), .IN4(n3361), .Q(
        n3198) );
  AO22X1 U2322 ( .IN1(n3561), .IN2(n3364), .IN3(elem30[3]), .IN4(n3361), .Q(
        n3199) );
  AO22X1 U2323 ( .IN1(n3564), .IN2(n3364), .IN3(elem30[4]), .IN4(n3361), .Q(
        n3200) );
  AO22X1 U2324 ( .IN1(n3567), .IN2(n3365), .IN3(elem30[5]), .IN4(n3361), .Q(
        n3201) );
  AO22X1 U2325 ( .IN1(n3570), .IN2(n3365), .IN3(elem30[6]), .IN4(n3361), .Q(
        n3202) );
  AO22X1 U2326 ( .IN1(n3573), .IN2(n3365), .IN3(elem30[7]), .IN4(n3361), .Q(
        n3203) );
  AO22X1 U2327 ( .IN1(n3576), .IN2(n3365), .IN3(elem30[8]), .IN4(n3361), .Q(
        n3204) );
  AO22X1 U2328 ( .IN1(n3579), .IN2(n3365), .IN3(elem30[9]), .IN4(n3361), .Q(
        n3205) );
  AO22X1 U2329 ( .IN1(n3582), .IN2(n3365), .IN3(elem30[10]), .IN4(n3361), .Q(
        n3206) );
  AO22X1 U2330 ( .IN1(n3585), .IN2(n3365), .IN3(elem30[11]), .IN4(n3361), .Q(
        n3207) );
  AND2X1 U2331 ( .IN1(n2230), .IN2(n2249), .Q(n2265) );
  AND2X1 U2332 ( .IN1(wr_en), .IN2(wr_addr[4]), .Q(n2230) );
  OR2X1 U2 ( .IN1(n993), .IN2(n994), .Q(rd_dataA[1]) );
  NAND4X0 U3 ( .IN1(n2009), .IN2(n2010), .IN3(n2011), .IN4(n2012), .QN(n993)
         );
  NAND4X0 U4 ( .IN1(n2002), .IN2(n2003), .IN3(n2004), .IN4(n2005), .QN(n994)
         );
  INVX0 U5 ( .INP(n2243), .ZN(n3298) );
  INVX0 U6 ( .INP(n2250), .ZN(n3278) );
  INVX0 U7 ( .INP(n2255), .ZN(n2000) );
  INVX0 U8 ( .INP(n2243), .ZN(n3299) );
  INVX0 U9 ( .INP(n2243), .ZN(n3300) );
  INVX0 U10 ( .INP(n2250), .ZN(n3279) );
  INVX0 U11 ( .INP(n2250), .ZN(n3280) );
  INVX0 U12 ( .INP(n2255), .ZN(n2001) );
  INVX0 U13 ( .INP(n2255), .ZN(n3260) );
  INVX0 U14 ( .INP(n2231), .ZN(n3338) );
  INVX0 U15 ( .INP(n2237), .ZN(n3318) );
  INVX0 U16 ( .INP(n2260), .ZN(n1020) );
  INVX0 U17 ( .INP(n2260), .ZN(n1021) );
  INVX0 U18 ( .INP(n2220), .ZN(n3360) );
  INVX0 U19 ( .INP(n2220), .ZN(n3359) );
  INVX0 U20 ( .INP(n2264), .ZN(n1007) );
  INVX0 U21 ( .INP(n2264), .ZN(n1008) );
  INVX0 U22 ( .INP(n2264), .ZN(n1009) );
  INVX0 U23 ( .INP(n2220), .ZN(n3358) );
  INVX0 U24 ( .INP(n2231), .ZN(n3339) );
  INVX0 U25 ( .INP(n2231), .ZN(n3340) );
  INVX0 U26 ( .INP(n2237), .ZN(n3319) );
  INVX0 U27 ( .INP(n2237), .ZN(n3320) );
  NBUFFX2 U28 ( .INP(n1675), .Z(n3369) );
  NBUFFX2 U29 ( .INP(n1675), .Z(n3370) );
  NBUFFX2 U30 ( .INP(n1668), .Z(n3385) );
  NBUFFX2 U31 ( .INP(n1663), .Z(n3397) );
  NBUFFX2 U32 ( .INP(n1673), .Z(n3373) );
  NBUFFX2 U33 ( .INP(n1668), .Z(n3384) );
  NBUFFX2 U34 ( .INP(n1663), .Z(n3396) );
  NBUFFX2 U35 ( .INP(n1673), .Z(n3372) );
  NBUFFX2 U36 ( .INP(n1675), .Z(n3371) );
  NBUFFX2 U37 ( .INP(n1668), .Z(n3386) );
  NBUFFX2 U38 ( .INP(n1663), .Z(n3398) );
  NBUFFX2 U39 ( .INP(n1673), .Z(n3374) );
  NBUFFX2 U40 ( .INP(n1085), .Z(n3463) );
  NBUFFX2 U41 ( .INP(n1085), .Z(n3464) );
  NBUFFX2 U42 ( .INP(n1085), .Z(n3462) );
  NBUFFX2 U43 ( .INP(n1078), .Z(n3478) );
  NBUFFX2 U44 ( .INP(n1073), .Z(n3490) );
  NBUFFX2 U45 ( .INP(n1083), .Z(n3466) );
  NBUFFX2 U46 ( .INP(n1078), .Z(n3477) );
  NBUFFX2 U47 ( .INP(n1073), .Z(n3489) );
  NBUFFX2 U48 ( .INP(n1083), .Z(n3465) );
  NBUFFX2 U49 ( .INP(n1078), .Z(n3479) );
  NBUFFX2 U50 ( .INP(n1073), .Z(n3491) );
  NBUFFX2 U51 ( .INP(n1083), .Z(n3467) );
  NAND2X1 U52 ( .IN1(n2244), .IN2(n2221), .QN(n2243) );
  NAND2X1 U53 ( .IN1(n2251), .IN2(n2221), .QN(n2250) );
  NAND2X1 U54 ( .IN1(n2256), .IN2(n2221), .QN(n2255) );
  INVX0 U55 ( .INP(n2245), .ZN(n3293) );
  INVX0 U56 ( .INP(n2246), .ZN(n3288) );
  INVX0 U57 ( .INP(n2252), .ZN(n3273) );
  INVX0 U58 ( .INP(n2253), .ZN(n3268) );
  INVX0 U59 ( .INP(n2257), .ZN(n1034) );
  INVX0 U60 ( .INP(n2258), .ZN(n1029) );
  INVX0 U61 ( .INP(n2247), .ZN(n3283) );
  INVX0 U62 ( .INP(n2254), .ZN(n3263) );
  INVX0 U63 ( .INP(n2259), .ZN(n1024) );
  NAND2X1 U64 ( .IN1(n2261), .IN2(n2221), .QN(n2260) );
  INVX0 U65 ( .INP(n2245), .ZN(n3294) );
  INVX0 U66 ( .INP(n2245), .ZN(n3295) );
  INVX0 U67 ( .INP(n2246), .ZN(n3289) );
  INVX0 U68 ( .INP(n2246), .ZN(n3290) );
  INVX0 U69 ( .INP(n2252), .ZN(n3274) );
  INVX0 U70 ( .INP(n2252), .ZN(n3275) );
  INVX0 U71 ( .INP(n2253), .ZN(n3269) );
  INVX0 U72 ( .INP(n2253), .ZN(n3270) );
  INVX0 U73 ( .INP(n2257), .ZN(n1035) );
  INVX0 U74 ( .INP(n2257), .ZN(n1036) );
  INVX0 U75 ( .INP(n2258), .ZN(n1030) );
  INVX0 U76 ( .INP(n2258), .ZN(n1031) );
  INVX0 U77 ( .INP(n2247), .ZN(n3284) );
  INVX0 U78 ( .INP(n2247), .ZN(n3285) );
  INVX0 U79 ( .INP(n2254), .ZN(n3264) );
  INVX0 U80 ( .INP(n2254), .ZN(n3265) );
  INVX0 U81 ( .INP(n2259), .ZN(n1025) );
  INVX0 U82 ( .INP(n2259), .ZN(n1026) );
  NAND2X1 U83 ( .IN1(n2232), .IN2(n2221), .QN(n2231) );
  NAND2X1 U84 ( .IN1(n2238), .IN2(n2221), .QN(n2237) );
  NAND2X1 U85 ( .IN1(n2221), .IN2(n2265), .QN(n2264) );
  NAND2X1 U86 ( .IN1(n2221), .IN2(n2222), .QN(n2220) );
  INVX0 U87 ( .INP(n2266), .ZN(n1002) );
  INVX0 U88 ( .INP(n2223), .ZN(n3353) );
  INVX0 U89 ( .INP(n2233), .ZN(n3333) );
  INVX0 U90 ( .INP(n2234), .ZN(n3328) );
  INVX0 U91 ( .INP(n2239), .ZN(n3313) );
  INVX0 U92 ( .INP(n2240), .ZN(n3308) );
  INVX0 U93 ( .INP(n2235), .ZN(n3323) );
  INVX0 U94 ( .INP(n2241), .ZN(n3303) );
  INVX0 U95 ( .INP(n2262), .ZN(n1016) );
  INVX0 U96 ( .INP(n2262), .ZN(n1017) );
  INVX0 U97 ( .INP(n2263), .ZN(n1012) );
  INVX0 U98 ( .INP(n2263), .ZN(n1013) );
  INVX0 U99 ( .INP(n2219), .ZN(n3365) );
  INVX0 U100 ( .INP(n2219), .ZN(n3363) );
  INVX0 U101 ( .INP(n2219), .ZN(n3364) );
  INVX0 U102 ( .INP(n2225), .ZN(n3348) );
  INVX0 U103 ( .INP(n2225), .ZN(n3349) );
  INVX0 U104 ( .INP(n2225), .ZN(n3350) );
  INVX0 U105 ( .INP(n2267), .ZN(n997) );
  INVX0 U106 ( .INP(n2267), .ZN(n998) );
  INVX0 U107 ( .INP(n2267), .ZN(n999) );
  INVX0 U108 ( .INP(n2227), .ZN(n3343) );
  INVX0 U109 ( .INP(n2227), .ZN(n3344) );
  INVX0 U110 ( .INP(n2227), .ZN(n3345) );
  INVX0 U111 ( .INP(n2266), .ZN(n1003) );
  INVX0 U112 ( .INP(n2266), .ZN(n1004) );
  INVX0 U113 ( .INP(n2223), .ZN(n3354) );
  INVX0 U114 ( .INP(n2223), .ZN(n3355) );
  INVX0 U115 ( .INP(n2233), .ZN(n3334) );
  INVX0 U116 ( .INP(n2233), .ZN(n3335) );
  INVX0 U117 ( .INP(n2234), .ZN(n3329) );
  INVX0 U118 ( .INP(n2234), .ZN(n3330) );
  INVX0 U119 ( .INP(n2239), .ZN(n3314) );
  INVX0 U120 ( .INP(n2239), .ZN(n3315) );
  INVX0 U121 ( .INP(n2240), .ZN(n3309) );
  INVX0 U122 ( .INP(n2240), .ZN(n3310) );
  INVX0 U123 ( .INP(n2235), .ZN(n3324) );
  INVX0 U124 ( .INP(n2235), .ZN(n3325) );
  INVX0 U125 ( .INP(n2241), .ZN(n3304) );
  INVX0 U126 ( .INP(n2241), .ZN(n3305) );
  NBUFFX2 U127 ( .INP(n3736), .Z(n3659) );
  NBUFFX2 U128 ( .INP(n3736), .Z(n3660) );
  NBUFFX2 U129 ( .INP(n3736), .Z(n3661) );
  NBUFFX2 U130 ( .INP(n3736), .Z(n3662) );
  NBUFFX2 U131 ( .INP(n3736), .Z(n3663) );
  NBUFFX2 U132 ( .INP(n3736), .Z(n3664) );
  NBUFFX2 U133 ( .INP(n3736), .Z(n3665) );
  NBUFFX2 U134 ( .INP(n3736), .Z(n3666) );
  NBUFFX2 U135 ( .INP(n3736), .Z(n3667) );
  NBUFFX2 U136 ( .INP(n3736), .Z(n3668) );
  NBUFFX2 U137 ( .INP(n3736), .Z(n3669) );
  NBUFFX2 U138 ( .INP(n3736), .Z(n3670) );
  NBUFFX2 U139 ( .INP(n3735), .Z(n3671) );
  NBUFFX2 U140 ( .INP(n3735), .Z(n3672) );
  NBUFFX2 U141 ( .INP(n3735), .Z(n3673) );
  NBUFFX2 U142 ( .INP(n3735), .Z(n3674) );
  NBUFFX2 U143 ( .INP(n3735), .Z(n3675) );
  NBUFFX2 U144 ( .INP(n3735), .Z(n3676) );
  NBUFFX2 U145 ( .INP(n3735), .Z(n3677) );
  NBUFFX2 U146 ( .INP(n3735), .Z(n3678) );
  NBUFFX2 U147 ( .INP(n3735), .Z(n3679) );
  NBUFFX2 U148 ( .INP(n3735), .Z(n3680) );
  NBUFFX2 U149 ( .INP(n3735), .Z(n3681) );
  NBUFFX2 U150 ( .INP(n3735), .Z(n3682) );
  NBUFFX2 U151 ( .INP(n3734), .Z(n3683) );
  NBUFFX2 U152 ( .INP(n3734), .Z(n3684) );
  NBUFFX2 U153 ( .INP(n3734), .Z(n3685) );
  NBUFFX2 U154 ( .INP(n3734), .Z(n3686) );
  NBUFFX2 U155 ( .INP(n3734), .Z(n3687) );
  NBUFFX2 U156 ( .INP(n3734), .Z(n3688) );
  NBUFFX2 U157 ( .INP(n3734), .Z(n3689) );
  NBUFFX2 U158 ( .INP(n3734), .Z(n3690) );
  NBUFFX2 U159 ( .INP(n3734), .Z(n3691) );
  NBUFFX2 U160 ( .INP(n3734), .Z(n3692) );
  NBUFFX2 U161 ( .INP(n3734), .Z(n3693) );
  NBUFFX2 U162 ( .INP(n3734), .Z(n3694) );
  NBUFFX2 U163 ( .INP(n3733), .Z(n3695) );
  NBUFFX2 U1108 ( .INP(n3733), .Z(n3696) );
  NBUFFX2 U1109 ( .INP(n3733), .Z(n3697) );
  NBUFFX2 U1117 ( .INP(n3733), .Z(n3698) );
  NBUFFX2 U2333 ( .INP(n3733), .Z(n3699) );
  NBUFFX2 U2334 ( .INP(n3733), .Z(n3700) );
  NBUFFX2 U2335 ( .INP(n3733), .Z(n3701) );
  NBUFFX2 U2336 ( .INP(n3733), .Z(n3702) );
  NBUFFX2 U2337 ( .INP(n3733), .Z(n3703) );
  NBUFFX2 U2338 ( .INP(n3733), .Z(n3704) );
  NBUFFX2 U2339 ( .INP(n3733), .Z(n3705) );
  NBUFFX2 U2340 ( .INP(n3733), .Z(n3706) );
  NBUFFX2 U2341 ( .INP(n3732), .Z(n3707) );
  NBUFFX2 U2342 ( .INP(n3732), .Z(n3708) );
  NBUFFX2 U2343 ( .INP(n3732), .Z(n3709) );
  NBUFFX2 U2344 ( .INP(n3732), .Z(n3710) );
  NBUFFX2 U2345 ( .INP(n3732), .Z(n3711) );
  NBUFFX2 U2346 ( .INP(n3732), .Z(n3712) );
  NBUFFX2 U2347 ( .INP(n3732), .Z(n3713) );
  NBUFFX2 U2348 ( .INP(n3732), .Z(n3714) );
  NBUFFX2 U2349 ( .INP(n3732), .Z(n3715) );
  NBUFFX2 U2350 ( .INP(n3732), .Z(n3716) );
  NBUFFX2 U2351 ( .INP(n3732), .Z(n3717) );
  NBUFFX2 U2352 ( .INP(n3732), .Z(n3718) );
  NBUFFX2 U2353 ( .INP(n3731), .Z(n3719) );
  NBUFFX2 U2354 ( .INP(n3731), .Z(n3720) );
  NBUFFX2 U2355 ( .INP(n3731), .Z(n3721) );
  NBUFFX2 U2356 ( .INP(n3731), .Z(n3722) );
  NBUFFX2 U2357 ( .INP(n3731), .Z(n3723) );
  NBUFFX2 U2358 ( .INP(n3731), .Z(n3724) );
  NBUFFX2 U2359 ( .INP(n3731), .Z(n3725) );
  NBUFFX2 U2360 ( .INP(n3731), .Z(n3726) );
  NBUFFX2 U2361 ( .INP(n3731), .Z(n3727) );
  NBUFFX2 U2362 ( .INP(n3731), .Z(n3728) );
  NBUFFX2 U2363 ( .INP(n3731), .Z(n3729) );
  NBUFFX2 U2364 ( .INP(n3737), .Z(n3648) );
  NBUFFX2 U2365 ( .INP(n3737), .Z(n3649) );
  NBUFFX2 U2366 ( .INP(n3737), .Z(n3650) );
  NBUFFX2 U2367 ( .INP(n3737), .Z(n3651) );
  NBUFFX2 U2368 ( .INP(n3737), .Z(n3652) );
  NBUFFX2 U2369 ( .INP(n3737), .Z(n3653) );
  NBUFFX2 U2370 ( .INP(n3737), .Z(n3654) );
  NBUFFX2 U2371 ( .INP(n3737), .Z(n3655) );
  NBUFFX2 U2372 ( .INP(n3737), .Z(n3656) );
  NBUFFX2 U2373 ( .INP(n3737), .Z(n3657) );
  NBUFFX2 U2374 ( .INP(n3737), .Z(n3658) );
  NBUFFX2 U2375 ( .INP(n3731), .Z(n3730) );
  NBUFFX2 U2376 ( .INP(n1670), .Z(n3382) );
  NBUFFX2 U2377 ( .INP(n1670), .Z(n3381) );
  NBUFFX2 U2378 ( .INP(n1665), .Z(n3393) );
  NBUFFX2 U2379 ( .INP(n1660), .Z(n3405) );
  NBUFFX2 U2380 ( .INP(n1665), .Z(n3394) );
  NBUFFX2 U2381 ( .INP(n1660), .Z(n3406) );
  NBUFFX2 U2382 ( .INP(n1638), .Z(n3451) );
  NBUFFX2 U2383 ( .INP(n1648), .Z(n3427) );
  NBUFFX2 U2384 ( .INP(n1643), .Z(n3439) );
  NBUFFX2 U2385 ( .INP(n1648), .Z(n3426) );
  NBUFFX2 U2386 ( .INP(n1643), .Z(n3438) );
  NBUFFX2 U2387 ( .INP(n1638), .Z(n3450) );
  NBUFFX2 U2388 ( .INP(n1650), .Z(n3421) );
  NBUFFX2 U2389 ( .INP(n1650), .Z(n3420) );
  NBUFFX2 U2390 ( .INP(n1666), .Z(n3391) );
  NBUFFX2 U2391 ( .INP(n1676), .Z(n3367) );
  NBUFFX2 U2392 ( .INP(n1671), .Z(n3379) );
  NBUFFX2 U2393 ( .INP(n1671), .Z(n3378) );
  NBUFFX2 U2394 ( .INP(n1666), .Z(n3390) );
  NBUFFX2 U2395 ( .INP(n1676), .Z(n3366) );
  NBUFFX2 U2396 ( .INP(n1661), .Z(n3403) );
  NBUFFX2 U2397 ( .INP(n1639), .Z(n3448) );
  NBUFFX2 U2398 ( .INP(n1661), .Z(n3402) );
  NBUFFX2 U2399 ( .INP(n1649), .Z(n3424) );
  NBUFFX2 U2400 ( .INP(n1644), .Z(n3436) );
  NBUFFX2 U2401 ( .INP(n1649), .Z(n3423) );
  NBUFFX2 U2402 ( .INP(n1644), .Z(n3435) );
  NBUFFX2 U2403 ( .INP(n1658), .Z(n3409) );
  NBUFFX2 U2404 ( .INP(n1658), .Z(n3408) );
  NBUFFX2 U2405 ( .INP(n1646), .Z(n3430) );
  NBUFFX2 U2406 ( .INP(n1641), .Z(n3442) );
  NBUFFX2 U2407 ( .INP(n1636), .Z(n3454) );
  NBUFFX2 U2408 ( .INP(n1646), .Z(n3429) );
  NBUFFX2 U2409 ( .INP(n1641), .Z(n3441) );
  NBUFFX2 U2410 ( .INP(n1636), .Z(n3453) );
  NBUFFX2 U2411 ( .INP(n1652), .Z(n3415) );
  NBUFFX2 U2412 ( .INP(n1652), .Z(n3414) );
  NBUFFX2 U2413 ( .INP(n1667), .Z(n3388) );
  NBUFFX2 U2414 ( .INP(n1662), .Z(n3400) );
  NBUFFX2 U2415 ( .INP(n1672), .Z(n3376) );
  NBUFFX2 U2416 ( .INP(n1657), .Z(n3412) );
  NBUFFX2 U2417 ( .INP(n1667), .Z(n3387) );
  NBUFFX2 U2418 ( .INP(n1662), .Z(n3399) );
  NBUFFX2 U2419 ( .INP(n1672), .Z(n3375) );
  NBUFFX2 U2420 ( .INP(n1657), .Z(n3411) );
  NBUFFX2 U2421 ( .INP(n1645), .Z(n3433) );
  NBUFFX2 U2422 ( .INP(n1640), .Z(n3445) );
  NBUFFX2 U2423 ( .INP(n1635), .Z(n3457) );
  NBUFFX2 U2424 ( .INP(n1645), .Z(n3432) );
  NBUFFX2 U2425 ( .INP(n1640), .Z(n3444) );
  NBUFFX2 U2426 ( .INP(n1635), .Z(n3456) );
  NBUFFX2 U2427 ( .INP(n1651), .Z(n3418) );
  NBUFFX2 U2428 ( .INP(n1651), .Z(n3417) );
  NBUFFX2 U2429 ( .INP(n1670), .Z(n3383) );
  NBUFFX2 U2430 ( .INP(n1665), .Z(n3395) );
  NBUFFX2 U2431 ( .INP(n1660), .Z(n3407) );
  NBUFFX2 U2432 ( .INP(n1648), .Z(n3428) );
  NBUFFX2 U2433 ( .INP(n1643), .Z(n3440) );
  NBUFFX2 U2434 ( .INP(n1638), .Z(n3452) );
  NBUFFX2 U2435 ( .INP(n1671), .Z(n3380) );
  NBUFFX2 U2436 ( .INP(n1666), .Z(n3392) );
  NBUFFX2 U2437 ( .INP(n1676), .Z(n3368) );
  NBUFFX2 U2438 ( .INP(n1661), .Z(n3404) );
  NBUFFX2 U2439 ( .INP(n1649), .Z(n3425) );
  NBUFFX2 U2440 ( .INP(n1644), .Z(n3437) );
  NAND2X1 U2441 ( .IN1(n2205), .IN2(n2212), .QN(n1675) );
  NAND2X1 U2442 ( .IN1(n2203), .IN2(n2212), .QN(n1668) );
  NAND2X1 U2443 ( .IN1(n2200), .IN2(n2212), .QN(n1663) );
  NAND2X1 U2444 ( .IN1(n2204), .IN2(n2212), .QN(n1673) );
  NBUFFX2 U2445 ( .INP(n1639), .Z(n3447) );
  NBUFFX2 U2446 ( .INP(n1650), .Z(n3422) );
  NBUFFX2 U2447 ( .INP(n1639), .Z(n3449) );
  NBUFFX2 U2448 ( .INP(n1658), .Z(n3410) );
  NBUFFX2 U2449 ( .INP(n1646), .Z(n3431) );
  NBUFFX2 U2450 ( .INP(n1641), .Z(n3443) );
  NBUFFX2 U2451 ( .INP(n1636), .Z(n3455) );
  NBUFFX2 U2452 ( .INP(n1652), .Z(n3416) );
  NBUFFX2 U2453 ( .INP(n1667), .Z(n3389) );
  NBUFFX2 U2454 ( .INP(n1662), .Z(n3401) );
  NBUFFX2 U2455 ( .INP(n1672), .Z(n3377) );
  NBUFFX2 U2456 ( .INP(n1657), .Z(n3413) );
  NBUFFX2 U2457 ( .INP(n1645), .Z(n3434) );
  NBUFFX2 U2458 ( .INP(n1640), .Z(n3446) );
  NBUFFX2 U2459 ( .INP(n1635), .Z(n3458) );
  NBUFFX2 U2460 ( .INP(n1651), .Z(n3419) );
  NBUFFX2 U2461 ( .INP(n1080), .Z(n3475) );
  NBUFFX2 U2462 ( .INP(n1075), .Z(n3487) );
  NBUFFX2 U2463 ( .INP(n1070), .Z(n3499) );
  NBUFFX2 U2464 ( .INP(n1053), .Z(n3532) );
  NBUFFX2 U2465 ( .INP(n1058), .Z(n3520) );
  NBUFFX2 U2466 ( .INP(n1048), .Z(n3544) );
  NBUFFX2 U2467 ( .INP(n1054), .Z(n3529) );
  NBUFFX2 U2468 ( .INP(n1081), .Z(n3472) );
  NBUFFX2 U2469 ( .INP(n1076), .Z(n3484) );
  NBUFFX2 U2470 ( .INP(n1080), .Z(n3476) );
  NBUFFX2 U2471 ( .INP(n1075), .Z(n3488) );
  NBUFFX2 U2472 ( .INP(n1070), .Z(n3500) );
  NBUFFX2 U2473 ( .INP(n1053), .Z(n3533) );
  NBUFFX2 U2474 ( .INP(n1058), .Z(n3521) );
  NBUFFX2 U2475 ( .INP(n1048), .Z(n3545) );
  NBUFFX2 U2476 ( .INP(n1054), .Z(n3530) );
  NBUFFX2 U2477 ( .INP(n1059), .Z(n3518) );
  NBUFFX2 U2478 ( .INP(n1081), .Z(n3473) );
  NBUFFX2 U2479 ( .INP(n1076), .Z(n3485) );
  NAND2X1 U2480 ( .IN1(n1615), .IN2(n1622), .QN(n1085) );
  NBUFFX2 U2481 ( .INP(n1080), .Z(n3474) );
  NBUFFX2 U2482 ( .INP(n1075), .Z(n3486) );
  NBUFFX2 U2483 ( .INP(n1070), .Z(n3498) );
  NBUFFX2 U2484 ( .INP(n1053), .Z(n3531) );
  NBUFFX2 U2485 ( .INP(n1058), .Z(n3519) );
  NBUFFX2 U2486 ( .INP(n1048), .Z(n3543) );
  NBUFFX2 U2487 ( .INP(n1071), .Z(n3496) );
  NBUFFX2 U2488 ( .INP(n1071), .Z(n3495) );
  NBUFFX2 U2489 ( .INP(n1059), .Z(n3517) );
  NBUFFX2 U2490 ( .INP(n1049), .Z(n3541) );
  NBUFFX2 U2491 ( .INP(n1054), .Z(n3528) );
  NBUFFX2 U2492 ( .INP(n1059), .Z(n3516) );
  NBUFFX2 U2493 ( .INP(n1086), .Z(n3460) );
  NBUFFX2 U2494 ( .INP(n1081), .Z(n3471) );
  NBUFFX2 U2495 ( .INP(n1076), .Z(n3483) );
  NBUFFX2 U2496 ( .INP(n1086), .Z(n3459) );
  NBUFFX2 U2497 ( .INP(n1077), .Z(n3481) );
  NBUFFX2 U2498 ( .INP(n1072), .Z(n3493) );
  NBUFFX2 U2499 ( .INP(n1082), .Z(n3469) );
  NBUFFX2 U2500 ( .INP(n1067), .Z(n3505) );
  NBUFFX2 U2501 ( .INP(n1077), .Z(n3480) );
  NBUFFX2 U2502 ( .INP(n1072), .Z(n3492) );
  NBUFFX2 U2503 ( .INP(n1082), .Z(n3468) );
  NBUFFX2 U2504 ( .INP(n1067), .Z(n3504) );
  NBUFFX2 U2505 ( .INP(n1050), .Z(n3538) );
  NBUFFX2 U2506 ( .INP(n1055), .Z(n3526) );
  NBUFFX2 U2507 ( .INP(n1045), .Z(n3550) );
  NBUFFX2 U2508 ( .INP(n1050), .Z(n3537) );
  NBUFFX2 U2509 ( .INP(n1055), .Z(n3525) );
  NBUFFX2 U2510 ( .INP(n1045), .Z(n3549) );
  NBUFFX2 U2511 ( .INP(n1051), .Z(n3535) );
  NBUFFX2 U2512 ( .INP(n1056), .Z(n3523) );
  NBUFFX2 U2513 ( .INP(n1046), .Z(n3547) );
  NBUFFX2 U2514 ( .INP(n1051), .Z(n3534) );
  NBUFFX2 U2515 ( .INP(n1056), .Z(n3522) );
  NBUFFX2 U2516 ( .INP(n1046), .Z(n3546) );
  NBUFFX2 U2517 ( .INP(n1068), .Z(n3502) );
  NBUFFX2 U2518 ( .INP(n1068), .Z(n3501) );
  NBUFFX2 U2519 ( .INP(n1062), .Z(n3508) );
  NBUFFX2 U2520 ( .INP(n1062), .Z(n3507) );
  NBUFFX2 U2521 ( .INP(n1060), .Z(n3514) );
  NBUFFX2 U2522 ( .INP(n1060), .Z(n3513) );
  NBUFFX2 U2523 ( .INP(n1061), .Z(n3511) );
  NBUFFX2 U2524 ( .INP(n1061), .Z(n3510) );
  NBUFFX2 U2525 ( .INP(n1071), .Z(n3497) );
  NBUFFX2 U2526 ( .INP(n1049), .Z(n3542) );
  NBUFFX2 U2527 ( .INP(n1086), .Z(n3461) );
  NBUFFX2 U2528 ( .INP(n1050), .Z(n3539) );
  NBUFFX2 U2529 ( .INP(n1055), .Z(n3527) );
  NBUFFX2 U2530 ( .INP(n1045), .Z(n3551) );
  NBUFFX2 U2531 ( .INP(n1077), .Z(n3482) );
  NBUFFX2 U2532 ( .INP(n1072), .Z(n3494) );
  NBUFFX2 U2533 ( .INP(n1082), .Z(n3470) );
  NBUFFX2 U2534 ( .INP(n1067), .Z(n3506) );
  NBUFFX2 U2535 ( .INP(n1051), .Z(n3536) );
  NBUFFX2 U2536 ( .INP(n1056), .Z(n3524) );
  NBUFFX2 U2537 ( .INP(n1046), .Z(n3548) );
  NBUFFX2 U2538 ( .INP(n1068), .Z(n3503) );
  NBUFFX2 U2539 ( .INP(n1062), .Z(n3509) );
  NBUFFX2 U2540 ( .INP(n1060), .Z(n3515) );
  NBUFFX2 U2541 ( .INP(n1061), .Z(n3512) );
  NAND2X1 U2542 ( .IN1(n1613), .IN2(n1622), .QN(n1078) );
  NAND2X1 U2543 ( .IN1(n1610), .IN2(n1622), .QN(n1073) );
  NAND2X1 U2544 ( .IN1(n1614), .IN2(n1622), .QN(n1083) );
  NBUFFX2 U2545 ( .INP(n1049), .Z(n3540) );
  NAND2X1 U2546 ( .IN1(n2244), .IN2(n2226), .QN(n2246) );
  NAND2X1 U2547 ( .IN1(n2251), .IN2(n2226), .QN(n2253) );
  NAND2X1 U2548 ( .IN1(n2256), .IN2(n2226), .QN(n2258) );
  NAND2X1 U2549 ( .IN1(n2244), .IN2(n2224), .QN(n2245) );
  NAND2X1 U2550 ( .IN1(n2251), .IN2(n2224), .QN(n2252) );
  NAND2X1 U2551 ( .IN1(n2256), .IN2(n2224), .QN(n2257) );
  NAND2X1 U2552 ( .IN1(n2244), .IN2(n2228), .QN(n2247) );
  NAND2X1 U2553 ( .IN1(n2251), .IN2(n2228), .QN(n2254) );
  NAND2X1 U2554 ( .IN1(n2256), .IN2(n2228), .QN(n2259) );
  NAND2X1 U2555 ( .IN1(n2261), .IN2(n2226), .QN(n2263) );
  NAND2X1 U2556 ( .IN1(n2261), .IN2(n2224), .QN(n2262) );
  NOR2X0 U2557 ( .IN1(n3739), .IN2(n3740), .QN(n2221) );
  NAND2X1 U2558 ( .IN1(n2232), .IN2(n2226), .QN(n2234) );
  NAND2X1 U2559 ( .IN1(n2238), .IN2(n2226), .QN(n2240) );
  NAND2X1 U2560 ( .IN1(n2222), .IN2(n2224), .QN(n2223) );
  NAND2X1 U2561 ( .IN1(n2232), .IN2(n2224), .QN(n2233) );
  NAND2X1 U2562 ( .IN1(n2238), .IN2(n2224), .QN(n2239) );
  NAND2X1 U2563 ( .IN1(n2232), .IN2(n2228), .QN(n2235) );
  NAND2X1 U2564 ( .IN1(n2238), .IN2(n2228), .QN(n2241) );
  NAND2X1 U2565 ( .IN1(n2226), .IN2(n2222), .QN(n2225) );
  NAND2X1 U2566 ( .IN1(n2226), .IN2(n2265), .QN(n2267) );
  NAND2X1 U2567 ( .IN1(n2224), .IN2(n2265), .QN(n2219) );
  NAND2X1 U2568 ( .IN1(n2228), .IN2(n2222), .QN(n2227) );
  NAND2X1 U2569 ( .IN1(n2228), .IN2(n2265), .QN(n2266) );
  NOR2X0 U2570 ( .IN1(n3742), .IN2(n3741), .QN(n2249) );
  NBUFFX2 U2571 ( .INP(nrst), .Z(n3736) );
  NBUFFX2 U2572 ( .INP(nrst), .Z(n3735) );
  NBUFFX2 U2573 ( .INP(nrst), .Z(n3734) );
  NBUFFX2 U2574 ( .INP(nrst), .Z(n3733) );
  NBUFFX2 U2575 ( .INP(nrst), .Z(n3732) );
  NBUFFX2 U2576 ( .INP(nrst), .Z(n3731) );
  NBUFFX2 U2577 ( .INP(nrst), .Z(n3737) );
  NOR2X0 U2578 ( .IN1(n3743), .IN2(n3747), .QN(n2212) );
  NAND2X0 U2579 ( .IN1(n2202), .IN2(n2212), .QN(n1670) );
  NAND2X0 U2580 ( .IN1(n2199), .IN2(n2212), .QN(n1665) );
  NAND2X0 U2581 ( .IN1(n2195), .IN2(n2212), .QN(n1660) );
  NAND2X0 U2582 ( .IN1(n2197), .IN2(n2212), .QN(n1658) );
  NAND2X0 U2583 ( .IN1(n2199), .IN2(n2211), .QN(n1666) );
  NAND2X1 U2584 ( .IN1(n2205), .IN2(n2211), .QN(n1676) );
  NAND2X0 U2585 ( .IN1(n2202), .IN2(n2211), .QN(n1671) );
  NAND2X1 U2586 ( .IN1(n2203), .IN2(n2211), .QN(n1667) );
  NAND2X1 U2587 ( .IN1(n2200), .IN2(n2211), .QN(n1662) );
  NAND2X1 U2588 ( .IN1(n2204), .IN2(n2211), .QN(n1672) );
  NAND2X1 U2589 ( .IN1(n2197), .IN2(n2211), .QN(n1657) );
  NAND2X1 U2590 ( .IN1(n2211), .IN2(n2195), .QN(n1661) );
  NAND2X1 U2591 ( .IN1(n2196), .IN2(n2195), .QN(n1638) );
  NAND2X0 U2592 ( .IN1(n2196), .IN2(n2202), .QN(n1648) );
  NAND2X0 U2593 ( .IN1(n2196), .IN2(n2199), .QN(n1643) );
  NAND2X1 U2594 ( .IN1(n2196), .IN2(n2205), .QN(n1650) );
  NAND2X1 U2595 ( .IN1(n2196), .IN2(n2204), .QN(n1651) );
  NAND2X1 U2596 ( .IN1(n2196), .IN2(n2203), .QN(n1646) );
  NAND2X1 U2597 ( .IN1(n2196), .IN2(n2200), .QN(n1641) );
  NAND2X1 U2598 ( .IN1(n2196), .IN2(n2197), .QN(n1636) );
  NAND2X0 U2599 ( .IN1(n2194), .IN2(n2202), .QN(n1649) );
  NAND2X0 U2600 ( .IN1(n2194), .IN2(n2199), .QN(n1644) );
  NAND2X1 U2601 ( .IN1(n2194), .IN2(n2204), .QN(n1652) );
  NAND2X1 U2602 ( .IN1(n2194), .IN2(n2195), .QN(n1639) );
  NAND2X1 U2603 ( .IN1(n2194), .IN2(n2203), .QN(n1645) );
  NAND2X1 U2604 ( .IN1(n2194), .IN2(n2200), .QN(n1640) );
  NAND2X1 U2605 ( .IN1(n2194), .IN2(n2197), .QN(n1635) );
  NOR2X0 U2606 ( .IN1(n3748), .IN2(n3752), .QN(n1622) );
  NBUFFX2 U2607 ( .INP(wr_data[0]), .Z(n3552) );
  NBUFFX2 U2608 ( .INP(wr_data[0]), .Z(n3553) );
  NAND2X1 U2609 ( .IN1(n1612), .IN2(n1622), .QN(n1080) );
  NAND2X1 U2610 ( .IN1(n1609), .IN2(n1622), .QN(n1075) );
  NAND2X1 U2611 ( .IN1(n1605), .IN2(n1622), .QN(n1070) );
  NAND2X1 U2612 ( .IN1(n1612), .IN2(n1621), .QN(n1081) );
  NAND2X1 U2613 ( .IN1(n1609), .IN2(n1621), .QN(n1076) );
  NAND2X1 U2614 ( .IN1(n1606), .IN2(n1609), .QN(n1053) );
  NAND2X1 U2615 ( .IN1(n1606), .IN2(n1612), .QN(n1058) );
  NAND2X1 U2616 ( .IN1(n1606), .IN2(n1605), .QN(n1048) );
  NAND2X1 U2617 ( .IN1(n1604), .IN2(n1609), .QN(n1054) );
  NAND2X1 U2618 ( .IN1(n1604), .IN2(n1612), .QN(n1059) );
  NBUFFX2 U2619 ( .INP(wr_data[31]), .Z(n3645) );
  NBUFFX2 U2620 ( .INP(wr_data[31]), .Z(n3646) );
  NBUFFX2 U2621 ( .INP(wr_data[0]), .Z(n3554) );
  NAND2X1 U2622 ( .IN1(n1607), .IN2(n1622), .QN(n1068) );
  NAND2X1 U2623 ( .IN1(n1615), .IN2(n1621), .QN(n1086) );
  NAND2X1 U2624 ( .IN1(n1613), .IN2(n1621), .QN(n1077) );
  NAND2X1 U2625 ( .IN1(n1610), .IN2(n1621), .QN(n1072) );
  NAND2X1 U2626 ( .IN1(n1614), .IN2(n1621), .QN(n1082) );
  NAND2X1 U2627 ( .IN1(n1607), .IN2(n1621), .QN(n1067) );
  NAND2X1 U2628 ( .IN1(n1621), .IN2(n1605), .QN(n1071) );
  NAND2X1 U2629 ( .IN1(n1606), .IN2(n1610), .QN(n1051) );
  NAND2X1 U2630 ( .IN1(n1606), .IN2(n1613), .QN(n1056) );
  NAND2X1 U2631 ( .IN1(n1606), .IN2(n1607), .QN(n1046) );
  NAND2X1 U2632 ( .IN1(n1606), .IN2(n1614), .QN(n1061) );
  NAND2X1 U2633 ( .IN1(n1606), .IN2(n1615), .QN(n1060) );
  NAND2X1 U2634 ( .IN1(n1604), .IN2(n1605), .QN(n1049) );
  NAND2X1 U2635 ( .IN1(n1604), .IN2(n1610), .QN(n1050) );
  NAND2X1 U2636 ( .IN1(n1604), .IN2(n1613), .QN(n1055) );
  NAND2X1 U2637 ( .IN1(n1604), .IN2(n1607), .QN(n1045) );
  NAND2X1 U2638 ( .IN1(n1604), .IN2(n1614), .QN(n1062) );
  NBUFFX2 U2639 ( .INP(wr_data[28]), .Z(n3636) );
  NBUFFX2 U2640 ( .INP(wr_data[29]), .Z(n3639) );
  NBUFFX2 U2641 ( .INP(wr_data[30]), .Z(n3642) );
  NBUFFX2 U2642 ( .INP(wr_data[28]), .Z(n3637) );
  NBUFFX2 U2643 ( .INP(wr_data[29]), .Z(n3640) );
  NBUFFX2 U2644 ( .INP(wr_data[30]), .Z(n3643) );
  NBUFFX2 U2645 ( .INP(wr_data[29]), .Z(n3641) );
  NBUFFX2 U2646 ( .INP(wr_data[30]), .Z(n3644) );
  NBUFFX2 U2647 ( .INP(wr_data[31]), .Z(n3647) );
  NBUFFX2 U2648 ( .INP(wr_data[24]), .Z(n3624) );
  NBUFFX2 U2649 ( .INP(wr_data[25]), .Z(n3627) );
  NBUFFX2 U2650 ( .INP(wr_data[26]), .Z(n3630) );
  NBUFFX2 U2651 ( .INP(wr_data[27]), .Z(n3633) );
  NBUFFX2 U2652 ( .INP(wr_data[24]), .Z(n3625) );
  NBUFFX2 U2653 ( .INP(wr_data[25]), .Z(n3628) );
  NBUFFX2 U2654 ( .INP(wr_data[26]), .Z(n3631) );
  NBUFFX2 U2655 ( .INP(wr_data[27]), .Z(n3634) );
  NBUFFX2 U2656 ( .INP(wr_data[25]), .Z(n3629) );
  NBUFFX2 U2657 ( .INP(wr_data[26]), .Z(n3632) );
  NBUFFX2 U2658 ( .INP(wr_data[27]), .Z(n3635) );
  NBUFFX2 U2659 ( .INP(wr_data[28]), .Z(n3638) );
  NBUFFX2 U2660 ( .INP(wr_data[20]), .Z(n3612) );
  NBUFFX2 U2661 ( .INP(wr_data[21]), .Z(n3615) );
  NBUFFX2 U2662 ( .INP(wr_data[22]), .Z(n3618) );
  NBUFFX2 U2663 ( .INP(wr_data[23]), .Z(n3621) );
  NBUFFX2 U2664 ( .INP(wr_data[20]), .Z(n3613) );
  NBUFFX2 U2665 ( .INP(wr_data[21]), .Z(n3616) );
  NBUFFX2 U2666 ( .INP(wr_data[22]), .Z(n3619) );
  NBUFFX2 U2667 ( .INP(wr_data[23]), .Z(n3622) );
  NBUFFX2 U2668 ( .INP(wr_data[21]), .Z(n3617) );
  NBUFFX2 U2669 ( .INP(wr_data[22]), .Z(n3620) );
  NBUFFX2 U2670 ( .INP(wr_data[23]), .Z(n3623) );
  NBUFFX2 U2671 ( .INP(wr_data[24]), .Z(n3626) );
  NBUFFX2 U2672 ( .INP(wr_data[17]), .Z(n3603) );
  NBUFFX2 U2673 ( .INP(wr_data[18]), .Z(n3606) );
  NBUFFX2 U2674 ( .INP(wr_data[19]), .Z(n3609) );
  NBUFFX2 U2675 ( .INP(wr_data[17]), .Z(n3604) );
  NBUFFX2 U2676 ( .INP(wr_data[18]), .Z(n3607) );
  NBUFFX2 U2677 ( .INP(wr_data[19]), .Z(n3610) );
  NBUFFX2 U2678 ( .INP(wr_data[18]), .Z(n3608) );
  NBUFFX2 U2679 ( .INP(wr_data[19]), .Z(n3611) );
  NBUFFX2 U2680 ( .INP(wr_data[20]), .Z(n3614) );
  NBUFFX2 U2681 ( .INP(wr_data[14]), .Z(n3594) );
  NBUFFX2 U2682 ( .INP(wr_data[15]), .Z(n3597) );
  NBUFFX2 U2683 ( .INP(wr_data[16]), .Z(n3600) );
  NBUFFX2 U2684 ( .INP(wr_data[13]), .Z(n3591) );
  NBUFFX2 U2685 ( .INP(wr_data[14]), .Z(n3595) );
  NBUFFX2 U2686 ( .INP(wr_data[15]), .Z(n3598) );
  NBUFFX2 U2687 ( .INP(wr_data[16]), .Z(n3601) );
  NBUFFX2 U2688 ( .INP(wr_data[13]), .Z(n3592) );
  NBUFFX2 U2689 ( .INP(wr_data[14]), .Z(n3596) );
  NBUFFX2 U2690 ( .INP(wr_data[15]), .Z(n3599) );
  NBUFFX2 U2691 ( .INP(wr_data[16]), .Z(n3602) );
  NBUFFX2 U2692 ( .INP(wr_data[17]), .Z(n3605) );
  NBUFFX2 U2693 ( .INP(wr_data[9]), .Z(n3579) );
  NBUFFX2 U2694 ( .INP(wr_data[10]), .Z(n3582) );
  NBUFFX2 U2695 ( .INP(wr_data[11]), .Z(n3585) );
  NBUFFX2 U2696 ( .INP(wr_data[12]), .Z(n3588) );
  NBUFFX2 U2697 ( .INP(wr_data[9]), .Z(n3580) );
  NBUFFX2 U2698 ( .INP(wr_data[12]), .Z(n3589) );
  NBUFFX2 U2699 ( .INP(wr_data[10]), .Z(n3583) );
  NBUFFX2 U2700 ( .INP(wr_data[11]), .Z(n3586) );
  NBUFFX2 U2701 ( .INP(wr_data[10]), .Z(n3584) );
  NBUFFX2 U2702 ( .INP(wr_data[11]), .Z(n3587) );
  NBUFFX2 U2703 ( .INP(wr_data[12]), .Z(n3590) );
  NBUFFX2 U2704 ( .INP(wr_data[13]), .Z(n3593) );
  NBUFFX2 U2705 ( .INP(wr_data[5]), .Z(n3567) );
  NBUFFX2 U2706 ( .INP(wr_data[6]), .Z(n3570) );
  NBUFFX2 U2707 ( .INP(wr_data[7]), .Z(n3573) );
  NBUFFX2 U2708 ( .INP(wr_data[8]), .Z(n3576) );
  NBUFFX2 U2709 ( .INP(wr_data[5]), .Z(n3568) );
  NBUFFX2 U2710 ( .INP(wr_data[6]), .Z(n3571) );
  NBUFFX2 U2711 ( .INP(wr_data[7]), .Z(n3574) );
  NBUFFX2 U2712 ( .INP(wr_data[8]), .Z(n3577) );
  NBUFFX2 U2713 ( .INP(wr_data[6]), .Z(n3572) );
  NBUFFX2 U2714 ( .INP(wr_data[7]), .Z(n3575) );
  NBUFFX2 U2715 ( .INP(wr_data[8]), .Z(n3578) );
  NBUFFX2 U2716 ( .INP(wr_data[9]), .Z(n3581) );
  NOR2X0 U2717 ( .IN1(n3738), .IN2(wr_addr[4]), .QN(n2248) );
  INVX0 U2718 ( .INP(wr_en), .ZN(n3738) );
  NBUFFX2 U2719 ( .INP(wr_data[2]), .Z(n3558) );
  NBUFFX2 U2720 ( .INP(wr_data[3]), .Z(n3561) );
  NBUFFX2 U2721 ( .INP(wr_data[4]), .Z(n3564) );
  NBUFFX2 U2722 ( .INP(wr_data[2]), .Z(n3559) );
  NBUFFX2 U2723 ( .INP(wr_data[3]), .Z(n3562) );
  NBUFFX2 U2724 ( .INP(wr_data[4]), .Z(n3565) );
  NBUFFX2 U2725 ( .INP(wr_data[3]), .Z(n3563) );
  NBUFFX2 U2726 ( .INP(wr_data[4]), .Z(n3566) );
  NBUFFX2 U2727 ( .INP(wr_data[5]), .Z(n3569) );
  NOR2X0 U2728 ( .IN1(n3739), .IN2(wr_addr[1]), .QN(n2226) );
  NOR2X0 U2729 ( .IN1(n3740), .IN2(wr_addr[0]), .QN(n2224) );
  NOR2X0 U2730 ( .IN1(wr_addr[0]), .IN2(wr_addr[1]), .QN(n2228) );
  NBUFFX2 U2731 ( .INP(wr_data[1]), .Z(n3555) );
  NBUFFX2 U2732 ( .INP(wr_data[1]), .Z(n3556) );
  INVX0 U2733 ( .INP(wr_addr[1]), .ZN(n3740) );
  INVX0 U2734 ( .INP(wr_addr[3]), .ZN(n3742) );
  NBUFFX2 U2735 ( .INP(wr_data[1]), .Z(n3557) );
  NBUFFX2 U2736 ( .INP(wr_data[2]), .Z(n3560) );
  INVX0 U2737 ( .INP(wr_addr[2]), .ZN(n3741) );
  INVX0 U2738 ( .INP(wr_addr[0]), .ZN(n3739) );
  NOR2X0 U2739 ( .IN1(n3741), .IN2(wr_addr[3]), .QN(n2236) );
  NOR2X0 U2740 ( .IN1(wr_addr[2]), .IN2(wr_addr[3]), .QN(n2242) );
  NOR2X0 U2741 ( .IN1(n3742), .IN2(wr_addr[2]), .QN(n2229) );
  NOR2X0 U2742 ( .IN1(n3743), .IN2(rd_addrA[0]), .QN(n2211) );
  NOR2X0 U2743 ( .IN1(n3747), .IN2(rd_addrA[4]), .QN(n2196) );
  NOR2X0 U2744 ( .IN1(rd_addrA[4]), .IN2(rd_addrA[0]), .QN(n2194) );
  INVX0 U2745 ( .INP(rd_addrA[0]), .ZN(n3747) );
  INVX0 U2746 ( .INP(rd_addrA[4]), .ZN(n3743) );
  NOR2X0 U2747 ( .IN1(n3745), .IN2(rd_addrA[1]), .QN(n2213) );
  NOR2X0 U2748 ( .IN1(n3744), .IN2(rd_addrA[2]), .QN(n2215) );
  NOR2X0 U2749 ( .IN1(n3746), .IN2(rd_addrA[3]), .QN(n2217) );
  INVX0 U2750 ( .INP(rd_addrA[3]), .ZN(n3744) );
  INVX0 U2751 ( .INP(rd_addrA[2]), .ZN(n3745) );
  INVX0 U2752 ( .INP(rd_addrA[1]), .ZN(n3746) );
  NOR2X0 U2753 ( .IN1(n3752), .IN2(rd_addrB[4]), .QN(n1606) );
  INVX0 U2754 ( .INP(rd_addrB[0]), .ZN(n3752) );
  INVX0 U2755 ( .INP(rd_addrB[4]), .ZN(n3748) );
  NOR2X0 U2756 ( .IN1(n3749), .IN2(rd_addrB[2]), .QN(n1625) );
  NOR2X0 U2757 ( .IN1(n3751), .IN2(rd_addrB[3]), .QN(n1627) );
  INVX0 U2758 ( .INP(rd_addrB[3]), .ZN(n3749) );
  INVX0 U2759 ( .INP(rd_addrB[1]), .ZN(n3751) );
  NOR2X0 U2760 ( .IN1(n3748), .IN2(rd_addrB[0]), .QN(n1621) );
  NOR2X0 U2761 ( .IN1(rd_addrB[4]), .IN2(rd_addrB[0]), .QN(n1604) );
  NOR2X0 U2762 ( .IN1(n3750), .IN2(rd_addrB[1]), .QN(n1623) );
  INVX0 U2763 ( .INP(rd_addrB[2]), .ZN(n3750) );
  INVX0 U2764 ( .INP(n998), .ZN(n995) );
  INVX0 U2765 ( .INP(n999), .ZN(n996) );
  INVX0 U2766 ( .INP(n1002), .ZN(n1000) );
  INVX0 U2767 ( .INP(n1002), .ZN(n1001) );
  INVX0 U2768 ( .INP(n1008), .ZN(n1005) );
  INVX0 U2769 ( .INP(n1009), .ZN(n1006) );
  INVX0 U2770 ( .INP(n1012), .ZN(n1010) );
  INVX0 U2771 ( .INP(n1013), .ZN(n1011) );
  INVX0 U2772 ( .INP(n1016), .ZN(n1014) );
  INVX0 U2773 ( .INP(n1017), .ZN(n1015) );
  INVX0 U2774 ( .INP(n1020), .ZN(n1018) );
  INVX0 U2775 ( .INP(n1021), .ZN(n1019) );
  INVX0 U2776 ( .INP(n1024), .ZN(n1022) );
  INVX0 U2777 ( .INP(n1024), .ZN(n1023) );
  INVX0 U2778 ( .INP(n1029), .ZN(n1027) );
  INVX0 U2779 ( .INP(n1029), .ZN(n1028) );
  INVX0 U2780 ( .INP(n1034), .ZN(n1032) );
  INVX0 U2781 ( .INP(n1034), .ZN(n1033) );
  INVX0 U2782 ( .INP(n2000), .ZN(n1037) );
  INVX0 U2783 ( .INP(n2000), .ZN(n1038) );
  INVX0 U2784 ( .INP(n3263), .ZN(n3261) );
  INVX0 U2785 ( .INP(n3263), .ZN(n3262) );
  INVX0 U2786 ( .INP(n3268), .ZN(n3266) );
  INVX0 U2787 ( .INP(n3268), .ZN(n3267) );
  INVX0 U2788 ( .INP(n3273), .ZN(n3271) );
  INVX0 U2789 ( .INP(n3273), .ZN(n3272) );
  INVX0 U2790 ( .INP(n3278), .ZN(n3276) );
  INVX0 U2791 ( .INP(n3278), .ZN(n3277) );
  INVX0 U2792 ( .INP(n3283), .ZN(n3281) );
  INVX0 U2793 ( .INP(n3283), .ZN(n3282) );
  INVX0 U2794 ( .INP(n3288), .ZN(n3286) );
  INVX0 U2795 ( .INP(n3288), .ZN(n3287) );
  INVX0 U2796 ( .INP(n3293), .ZN(n3291) );
  INVX0 U2797 ( .INP(n3293), .ZN(n3292) );
  INVX0 U2798 ( .INP(n3298), .ZN(n3296) );
  INVX0 U2799 ( .INP(n3298), .ZN(n3297) );
  INVX0 U2800 ( .INP(n3303), .ZN(n3301) );
  INVX0 U2801 ( .INP(n3303), .ZN(n3302) );
  INVX0 U2802 ( .INP(n3308), .ZN(n3306) );
  INVX0 U2803 ( .INP(n3308), .ZN(n3307) );
  INVX0 U2804 ( .INP(n3313), .ZN(n3311) );
  INVX0 U2805 ( .INP(n3313), .ZN(n3312) );
  INVX0 U2806 ( .INP(n3318), .ZN(n3316) );
  INVX0 U2807 ( .INP(n3318), .ZN(n3317) );
  INVX0 U2808 ( .INP(n3323), .ZN(n3321) );
  INVX0 U2809 ( .INP(n3323), .ZN(n3322) );
  INVX0 U2810 ( .INP(n3328), .ZN(n3326) );
  INVX0 U2811 ( .INP(n3328), .ZN(n3327) );
  INVX0 U2812 ( .INP(n3333), .ZN(n3331) );
  INVX0 U2813 ( .INP(n3333), .ZN(n3332) );
  INVX0 U2814 ( .INP(n3338), .ZN(n3336) );
  INVX0 U2815 ( .INP(n3338), .ZN(n3337) );
  INVX0 U2816 ( .INP(n3344), .ZN(n3341) );
  INVX0 U2817 ( .INP(n3345), .ZN(n3342) );
  INVX0 U2818 ( .INP(n3349), .ZN(n3346) );
  INVX0 U2819 ( .INP(n3350), .ZN(n3347) );
  INVX0 U2820 ( .INP(n3353), .ZN(n3351) );
  INVX0 U2821 ( .INP(n3353), .ZN(n3352) );
  INVX0 U2822 ( .INP(n3359), .ZN(n3356) );
  INVX0 U2823 ( .INP(n3358), .ZN(n3357) );
  INVX0 U2824 ( .INP(n3363), .ZN(n3361) );
  INVX0 U2825 ( .INP(n3364), .ZN(n3362) );
endmodule


module single_cycle_mips_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_31 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry[31]), .Q(SUM[31]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module single_cycle_mips_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [31:1] carry;

  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n15), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(A[21]), .IN2(n2), .Q(n1) );
  AND2X1 U2 ( .IN1(A[20]), .IN2(n4), .Q(n2) );
  AND2X1 U3 ( .IN1(A[24]), .IN2(n5), .Q(n3) );
  AND2X1 U4 ( .IN1(A[19]), .IN2(n6), .Q(n4) );
  AND2X1 U5 ( .IN1(A[23]), .IN2(n7), .Q(n5) );
  NAND2X1 U6 ( .IN1(A[30]), .IN2(n12), .QN(n16) );
  AND2X1 U7 ( .IN1(A[18]), .IN2(n8), .Q(n6) );
  AND2X1 U8 ( .IN1(A[22]), .IN2(n1), .Q(n7) );
  AND2X1 U9 ( .IN1(A[17]), .IN2(n14), .Q(n8) );
  AND2X1 U10 ( .IN1(A[25]), .IN2(n3), .Q(n9) );
  AND2X1 U11 ( .IN1(A[28]), .IN2(n11), .Q(n10) );
  AND2X1 U12 ( .IN1(A[27]), .IN2(n13), .Q(n11) );
  AND2X1 U13 ( .IN1(A[29]), .IN2(n10), .Q(n12) );
  AND2X1 U14 ( .IN1(A[26]), .IN2(n9), .Q(n13) );
  AND2X1 U15 ( .IN1(A[16]), .IN2(carry[16]), .Q(n14) );
  XNOR2X1 U16 ( .IN1(A[31]), .IN2(n16), .Q(SUM[31]) );
  AND2X1 U17 ( .IN1(A[0]), .IN2(B[0]), .Q(n15) );
  XOR2X1 U18 ( .IN1(A[30]), .IN2(n12), .Q(SUM[30]) );
  XOR2X1 U19 ( .IN1(A[29]), .IN2(n10), .Q(SUM[29]) );
  XOR2X1 U20 ( .IN1(A[28]), .IN2(n11), .Q(SUM[28]) );
  XOR2X1 U21 ( .IN1(A[27]), .IN2(n13), .Q(SUM[27]) );
  XOR2X1 U22 ( .IN1(A[26]), .IN2(n9), .Q(SUM[26]) );
  XOR2X1 U23 ( .IN1(A[25]), .IN2(n3), .Q(SUM[25]) );
  XOR2X1 U24 ( .IN1(A[24]), .IN2(n5), .Q(SUM[24]) );
  XOR2X1 U25 ( .IN1(A[23]), .IN2(n7), .Q(SUM[23]) );
  XOR2X1 U26 ( .IN1(A[22]), .IN2(n1), .Q(SUM[22]) );
  XOR2X1 U27 ( .IN1(A[21]), .IN2(n2), .Q(SUM[21]) );
  XOR2X1 U28 ( .IN1(A[20]), .IN2(n4), .Q(SUM[20]) );
  XOR2X1 U29 ( .IN1(A[19]), .IN2(n6), .Q(SUM[19]) );
  XOR2X1 U30 ( .IN1(A[18]), .IN2(n8), .Q(SUM[18]) );
  XOR2X1 U31 ( .IN1(A[17]), .IN2(n14), .Q(SUM[17]) );
  XOR2X1 U32 ( .IN1(A[16]), .IN2(carry[16]), .Q(SUM[16]) );
  XOR2X1 U33 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module single_cycle_mips_DW01_add_2 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_31 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry[31]), .Q(SUM[31]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module single_cycle_mips_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   \carry[31] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52;

  INVX0 U1 ( .INP(A[2]), .ZN(n14) );
  INVX0 U2 ( .INP(A[4]), .ZN(n12) );
  INVX0 U3 ( .INP(A[6]), .ZN(n10) );
  INVX0 U4 ( .INP(A[8]), .ZN(n8) );
  INVX0 U5 ( .INP(A[10]), .ZN(n6) );
  INVX0 U6 ( .INP(A[12]), .ZN(n4) );
  INVX0 U7 ( .INP(A[14]), .ZN(n2) );
  INVX0 U8 ( .INP(A[15]), .ZN(n1) );
  XNOR2X1 U9 ( .IN1(\carry[31] ), .IN2(A[31]), .Q(DIFF[31]) );
  INVX0 U10 ( .INP(A[1]), .ZN(n15) );
  INVX0 U11 ( .INP(A[3]), .ZN(n13) );
  INVX0 U12 ( .INP(A[5]), .ZN(n11) );
  INVX0 U13 ( .INP(A[7]), .ZN(n9) );
  INVX0 U14 ( .INP(A[9]), .ZN(n7) );
  INVX0 U15 ( .INP(A[11]), .ZN(n5) );
  INVX0 U16 ( .INP(A[13]), .ZN(n3) );
  INVX0 U17 ( .INP(B[0]), .ZN(n16) );
  NAND4X0 U18 ( .IN1(n17), .IN2(n18), .IN3(n19), .IN4(n20), .QN(\carry[31] )
         );
  NOR4X0 U19 ( .IN1(n21), .IN2(A[28]), .IN3(A[30]), .IN4(A[29]), .QN(n20) );
  OR2X1 U20 ( .IN1(A[27]), .IN2(A[26]), .Q(n21) );
  NOR4X0 U21 ( .IN1(A[25]), .IN2(A[24]), .IN3(A[23]), .IN4(A[22]), .QN(n19) );
  NOR4X0 U22 ( .IN1(A[21]), .IN2(A[20]), .IN3(A[19]), .IN4(A[18]), .QN(n18) );
  OA221X1 U23 ( .IN1(n22), .IN2(n1), .IN3(B[15]), .IN4(n23), .IN5(n24), .Q(n17) );
  NOR2X0 U24 ( .IN1(A[17]), .IN2(A[16]), .QN(n24) );
  AND2X1 U25 ( .IN1(n1), .IN2(n22), .Q(n23) );
  OA22X1 U26 ( .IN1(n25), .IN2(n2), .IN3(B[14]), .IN4(n26), .Q(n22) );
  AND2X1 U27 ( .IN1(n2), .IN2(n25), .Q(n26) );
  OA22X1 U28 ( .IN1(n27), .IN2(n3), .IN3(B[13]), .IN4(n28), .Q(n25) );
  AND2X1 U29 ( .IN1(n3), .IN2(n27), .Q(n28) );
  OA22X1 U30 ( .IN1(n29), .IN2(n4), .IN3(B[12]), .IN4(n30), .Q(n27) );
  AND2X1 U31 ( .IN1(n4), .IN2(n29), .Q(n30) );
  OA22X1 U32 ( .IN1(n31), .IN2(n5), .IN3(B[11]), .IN4(n32), .Q(n29) );
  AND2X1 U33 ( .IN1(n5), .IN2(n31), .Q(n32) );
  OA22X1 U34 ( .IN1(n33), .IN2(n6), .IN3(B[10]), .IN4(n34), .Q(n31) );
  AND2X1 U35 ( .IN1(n6), .IN2(n33), .Q(n34) );
  OA22X1 U36 ( .IN1(n35), .IN2(n7), .IN3(B[9]), .IN4(n36), .Q(n33) );
  AND2X1 U37 ( .IN1(n7), .IN2(n35), .Q(n36) );
  OA22X1 U38 ( .IN1(n37), .IN2(n8), .IN3(B[8]), .IN4(n38), .Q(n35) );
  AND2X1 U39 ( .IN1(n8), .IN2(n37), .Q(n38) );
  OA22X1 U40 ( .IN1(n39), .IN2(n9), .IN3(B[7]), .IN4(n40), .Q(n37) );
  AND2X1 U41 ( .IN1(n9), .IN2(n39), .Q(n40) );
  OA22X1 U42 ( .IN1(n41), .IN2(n10), .IN3(B[6]), .IN4(n42), .Q(n39) );
  AND2X1 U43 ( .IN1(n10), .IN2(n41), .Q(n42) );
  OA22X1 U44 ( .IN1(n43), .IN2(n11), .IN3(B[5]), .IN4(n44), .Q(n41) );
  AND2X1 U45 ( .IN1(n11), .IN2(n43), .Q(n44) );
  OA22X1 U46 ( .IN1(n45), .IN2(n12), .IN3(B[4]), .IN4(n46), .Q(n43) );
  AND2X1 U47 ( .IN1(n12), .IN2(n45), .Q(n46) );
  OA22X1 U48 ( .IN1(n47), .IN2(n13), .IN3(B[3]), .IN4(n48), .Q(n45) );
  AND2X1 U49 ( .IN1(n13), .IN2(n47), .Q(n48) );
  OA22X1 U50 ( .IN1(n49), .IN2(n14), .IN3(B[2]), .IN4(n50), .Q(n47) );
  AND2X1 U51 ( .IN1(n14), .IN2(n49), .Q(n50) );
  OA22X1 U52 ( .IN1(n51), .IN2(n15), .IN3(B[1]), .IN4(n52), .Q(n49) );
  AND2X1 U53 ( .IN1(n15), .IN2(n51), .Q(n52) );
  NOR2X0 U54 ( .IN1(n16), .IN2(A[0]), .QN(n51) );
endmodule


module single_cycle_mips_DW01_add_3 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  XOR3X1 U1_31 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry[31]), .Q(SUM[31]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module single_cycle_mips_DW01_add_4 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;
  assign SUM[1] = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  AND2X1 U1 ( .IN1(A[30]), .IN2(n24), .Q(n1) );
  INVX0 U2 ( .INP(A[2]), .ZN(SUM[2]) );
  AND2X1 U3 ( .IN1(A[4]), .IN2(n25), .Q(n2) );
  AND2X1 U4 ( .IN1(A[5]), .IN2(n2), .Q(n3) );
  AND2X1 U5 ( .IN1(A[6]), .IN2(n3), .Q(n4) );
  AND2X1 U6 ( .IN1(A[7]), .IN2(n4), .Q(n5) );
  AND2X1 U7 ( .IN1(A[8]), .IN2(n5), .Q(n6) );
  AND2X1 U8 ( .IN1(A[9]), .IN2(n6), .Q(n7) );
  AND2X1 U9 ( .IN1(A[10]), .IN2(n7), .Q(n8) );
  AND2X1 U10 ( .IN1(A[12]), .IN2(n26), .Q(n9) );
  AND2X1 U11 ( .IN1(A[13]), .IN2(n9), .Q(n10) );
  AND2X1 U12 ( .IN1(A[14]), .IN2(n10), .Q(n11) );
  AND2X1 U13 ( .IN1(A[16]), .IN2(n27), .Q(n12) );
  AND2X1 U14 ( .IN1(A[17]), .IN2(n12), .Q(n13) );
  AND2X1 U15 ( .IN1(A[18]), .IN2(n13), .Q(n14) );
  AND2X1 U16 ( .IN1(A[19]), .IN2(n14), .Q(n15) );
  AND2X1 U17 ( .IN1(A[20]), .IN2(n15), .Q(n16) );
  AND2X1 U18 ( .IN1(A[21]), .IN2(n16), .Q(n17) );
  AND2X1 U19 ( .IN1(A[22]), .IN2(n17), .Q(n18) );
  AND2X1 U20 ( .IN1(A[24]), .IN2(n28), .Q(n19) );
  AND2X1 U21 ( .IN1(A[25]), .IN2(n19), .Q(n20) );
  AND2X1 U22 ( .IN1(A[26]), .IN2(n20), .Q(n21) );
  AND2X1 U23 ( .IN1(A[27]), .IN2(n21), .Q(n22) );
  AND2X1 U24 ( .IN1(A[28]), .IN2(n22), .Q(n23) );
  AND2X1 U25 ( .IN1(A[29]), .IN2(n23), .Q(n24) );
  AND2X1 U26 ( .IN1(A[3]), .IN2(A[2]), .Q(n25) );
  AND2X1 U27 ( .IN1(A[11]), .IN2(n8), .Q(n26) );
  AND2X1 U28 ( .IN1(A[15]), .IN2(n11), .Q(n27) );
  AND2X1 U29 ( .IN1(A[23]), .IN2(n18), .Q(n28) );
  XOR2X1 U30 ( .IN1(A[31]), .IN2(n1), .Q(SUM[31]) );
  XOR2X1 U31 ( .IN1(A[30]), .IN2(n24), .Q(SUM[30]) );
  XOR2X1 U32 ( .IN1(A[29]), .IN2(n23), .Q(SUM[29]) );
  XOR2X1 U33 ( .IN1(A[28]), .IN2(n22), .Q(SUM[28]) );
  XOR2X1 U34 ( .IN1(A[27]), .IN2(n21), .Q(SUM[27]) );
  XOR2X1 U35 ( .IN1(A[26]), .IN2(n20), .Q(SUM[26]) );
  XOR2X1 U36 ( .IN1(A[25]), .IN2(n19), .Q(SUM[25]) );
  XOR2X1 U37 ( .IN1(A[24]), .IN2(n28), .Q(SUM[24]) );
  XOR2X1 U38 ( .IN1(A[23]), .IN2(n18), .Q(SUM[23]) );
  XOR2X1 U39 ( .IN1(A[22]), .IN2(n17), .Q(SUM[22]) );
  XOR2X1 U40 ( .IN1(A[21]), .IN2(n16), .Q(SUM[21]) );
  XOR2X1 U41 ( .IN1(A[20]), .IN2(n15), .Q(SUM[20]) );
  XOR2X1 U42 ( .IN1(A[19]), .IN2(n14), .Q(SUM[19]) );
  XOR2X1 U43 ( .IN1(A[18]), .IN2(n13), .Q(SUM[18]) );
  XOR2X1 U44 ( .IN1(A[17]), .IN2(n12), .Q(SUM[17]) );
  XOR2X1 U45 ( .IN1(A[16]), .IN2(n27), .Q(SUM[16]) );
  XOR2X1 U46 ( .IN1(A[15]), .IN2(n11), .Q(SUM[15]) );
  XOR2X1 U47 ( .IN1(A[14]), .IN2(n10), .Q(SUM[14]) );
  XOR2X1 U48 ( .IN1(A[13]), .IN2(n9), .Q(SUM[13]) );
  XOR2X1 U49 ( .IN1(A[12]), .IN2(n26), .Q(SUM[12]) );
  XOR2X1 U50 ( .IN1(A[11]), .IN2(n8), .Q(SUM[11]) );
  XOR2X1 U51 ( .IN1(A[10]), .IN2(n7), .Q(SUM[10]) );
  XOR2X1 U52 ( .IN1(A[9]), .IN2(n6), .Q(SUM[9]) );
  XOR2X1 U53 ( .IN1(A[8]), .IN2(n5), .Q(SUM[8]) );
  XOR2X1 U54 ( .IN1(A[7]), .IN2(n4), .Q(SUM[7]) );
  XOR2X1 U55 ( .IN1(A[6]), .IN2(n3), .Q(SUM[6]) );
  XOR2X1 U56 ( .IN1(A[5]), .IN2(n2), .Q(SUM[5]) );
  XOR2X1 U57 ( .IN1(A[4]), .IN2(n25), .Q(SUM[4]) );
  XOR2X1 U58 ( .IN1(A[3]), .IN2(A[2]), .Q(SUM[3]) );
endmodule


module single_cycle_mips_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [32:0] carry;

  FADDX1 U2_30 ( .A(A[30]), .B(n2), .CI(carry[30]), .CO(carry[31]), .S(
        DIFF[30]) );
  FADDX1 U2_29 ( .A(A[29]), .B(n2), .CI(carry[29]), .CO(carry[30]), .S(
        DIFF[29]) );
  FADDX1 U2_28 ( .A(A[28]), .B(n2), .CI(carry[28]), .CO(carry[29]), .S(
        DIFF[28]) );
  FADDX1 U2_27 ( .A(A[27]), .B(n2), .CI(carry[27]), .CO(carry[28]), .S(
        DIFF[27]) );
  FADDX1 U2_26 ( .A(A[26]), .B(n2), .CI(carry[26]), .CO(carry[27]), .S(
        DIFF[26]) );
  FADDX1 U2_25 ( .A(A[25]), .B(n2), .CI(carry[25]), .CO(carry[26]), .S(
        DIFF[25]) );
  FADDX1 U2_24 ( .A(A[24]), .B(n2), .CI(carry[24]), .CO(carry[25]), .S(
        DIFF[24]) );
  FADDX1 U2_23 ( .A(A[23]), .B(n2), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1 U2_22 ( .A(A[22]), .B(n2), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1 U2_21 ( .A(A[21]), .B(n2), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1 U2_20 ( .A(A[20]), .B(n2), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1 U2_19 ( .A(A[19]), .B(n2), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1 U2_18 ( .A(A[18]), .B(n2), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1 U2_17 ( .A(A[17]), .B(n2), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1 U2_16 ( .A(A[16]), .B(n2), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1 U2_15 ( .A(A[15]), .B(n2), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1 U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_31 ( .IN1(A[31]), .IN2(n2), .IN3(carry[31]), .Q(DIFF[31]) );
  INVX0 U1 ( .INP(B[3]), .ZN(n14) );
  INVX0 U2 ( .INP(B[4]), .ZN(n13) );
  INVX0 U3 ( .INP(B[5]), .ZN(n12) );
  INVX0 U4 ( .INP(B[2]), .ZN(n15) );
  INVX0 U5 ( .INP(B[9]), .ZN(n8) );
  INVX0 U6 ( .INP(B[8]), .ZN(n9) );
  INVX0 U7 ( .INP(B[7]), .ZN(n10) );
  INVX0 U8 ( .INP(B[6]), .ZN(n11) );
  INVX0 U9 ( .INP(B[1]), .ZN(n16) );
  NAND2X1 U10 ( .IN1(n1), .IN2(B[0]), .QN(carry[1]) );
  INVX0 U11 ( .INP(A[0]), .ZN(n1) );
  INVX0 U12 ( .INP(B[14]), .ZN(n3) );
  INVX0 U13 ( .INP(B[13]), .ZN(n4) );
  INVX0 U14 ( .INP(B[12]), .ZN(n5) );
  INVX0 U15 ( .INP(B[11]), .ZN(n6) );
  INVX0 U16 ( .INP(B[10]), .ZN(n7) );
  XOR2X1 U17 ( .IN1(B[0]), .IN2(A[0]), .Q(DIFF[0]) );
  INVX1 U18 ( .INP(B[31]), .ZN(n2) );
endmodule


module single_cycle_mips ( clk, rst_n, inst_addr, inst, data_addr, data_in, 
        data_out, data_wr );
  output [31:0] inst_addr;
  input [31:0] inst;
  output [31:0] data_addr;
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst_n;
  output data_wr;
  wire   N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36,
         N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50,
         N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64,
         N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78,
         N79, N80, N81, N82, N83, N84, N85, N86, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, wr_en, \diff_immed[31] , N191, N192,
         N193, N194, N195, N196, N197, N198, N199, N200, N201, N202, N203,
         N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, N214,
         N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N239, N240, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N378, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160;
  wire   [4:0] wr_addr;
  wire   [31:0] wr_data;
  wire   [31:0] rd_dataA;
  wire   [31:0] diff;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  DFFARX1 \pc_reg[0]  ( .D(N119), .CLK(clk), .RSTB(n144), .Q(inst_addr[0]) );
  DFFARX1 \pc_reg[1]  ( .D(N120), .CLK(clk), .RSTB(n144), .Q(inst_addr[1]) );
  DFFARX1 \pc_reg[2]  ( .D(N121), .CLK(clk), .RSTB(n144), .Q(inst_addr[2]) );
  DFFARX1 \pc_reg[3]  ( .D(N122), .CLK(clk), .RSTB(n144), .Q(inst_addr[3]) );
  DFFARX1 \pc_reg[4]  ( .D(N123), .CLK(clk), .RSTB(n144), .Q(inst_addr[4]) );
  DFFARX1 \pc_reg[5]  ( .D(N124), .CLK(clk), .RSTB(n144), .Q(inst_addr[5]) );
  DFFARX1 \pc_reg[6]  ( .D(N125), .CLK(clk), .RSTB(n144), .Q(inst_addr[6]) );
  DFFARX1 \pc_reg[7]  ( .D(N126), .CLK(clk), .RSTB(n144), .Q(inst_addr[7]) );
  DFFARX1 \pc_reg[8]  ( .D(N127), .CLK(clk), .RSTB(n144), .Q(inst_addr[8]) );
  DFFARX1 \pc_reg[9]  ( .D(N128), .CLK(clk), .RSTB(n144), .Q(inst_addr[9]) );
  DFFARX1 \pc_reg[10]  ( .D(N129), .CLK(clk), .RSTB(n144), .Q(inst_addr[10])
         );
  DFFARX1 \pc_reg[11]  ( .D(N130), .CLK(clk), .RSTB(n144), .Q(inst_addr[11])
         );
  DFFARX1 \pc_reg[12]  ( .D(N131), .CLK(clk), .RSTB(n144), .Q(inst_addr[12])
         );
  DFFARX1 \pc_reg[13]  ( .D(N132), .CLK(clk), .RSTB(n144), .Q(inst_addr[13])
         );
  DFFARX1 \pc_reg[14]  ( .D(N133), .CLK(clk), .RSTB(n144), .Q(inst_addr[14])
         );
  DFFARX1 \pc_reg[15]  ( .D(N134), .CLK(clk), .RSTB(n144), .Q(inst_addr[15])
         );
  DFFARX1 \pc_reg[16]  ( .D(N135), .CLK(clk), .RSTB(n144), .Q(inst_addr[16])
         );
  DFFARX1 \pc_reg[17]  ( .D(N136), .CLK(clk), .RSTB(n122), .Q(inst_addr[17])
         );
  DFFARX1 \pc_reg[18]  ( .D(N137), .CLK(clk), .RSTB(n122), .Q(inst_addr[18])
         );
  DFFARX1 \pc_reg[19]  ( .D(N138), .CLK(clk), .RSTB(n122), .Q(inst_addr[19])
         );
  DFFARX1 \pc_reg[20]  ( .D(N139), .CLK(clk), .RSTB(n122), .Q(inst_addr[20])
         );
  DFFARX1 \pc_reg[21]  ( .D(N140), .CLK(clk), .RSTB(n122), .Q(inst_addr[21])
         );
  DFFARX1 \pc_reg[22]  ( .D(N141), .CLK(clk), .RSTB(n122), .Q(inst_addr[22])
         );
  DFFARX1 \pc_reg[23]  ( .D(N142), .CLK(clk), .RSTB(n122), .Q(inst_addr[23])
         );
  DFFARX1 \pc_reg[24]  ( .D(N143), .CLK(clk), .RSTB(n122), .Q(inst_addr[24])
         );
  DFFARX1 \pc_reg[25]  ( .D(N144), .CLK(clk), .RSTB(n122), .Q(inst_addr[25])
         );
  DFFARX1 \pc_reg[26]  ( .D(N145), .CLK(clk), .RSTB(n122), .Q(inst_addr[26])
         );
  DFFARX1 \pc_reg[27]  ( .D(N146), .CLK(clk), .RSTB(n122), .Q(inst_addr[27])
         );
  DFFARX1 \pc_reg[28]  ( .D(N147), .CLK(clk), .RSTB(n122), .Q(inst_addr[28])
         );
  DFFARX1 \pc_reg[29]  ( .D(N148), .CLK(clk), .RSTB(n122), .Q(inst_addr[29])
         );
  DFFARX1 \pc_reg[30]  ( .D(N149), .CLK(clk), .RSTB(n122), .Q(inst_addr[30])
         );
  DFFARX1 \pc_reg[31]  ( .D(N150), .CLK(clk), .RSTB(n122), .Q(inst_addr[31])
         );
  OR4X1 U23 ( .IN1(n135), .IN2(n133), .IN3(n131), .IN4(n70), .Q(wr_en) );
  AO21X1 U24 ( .IN1(n71), .IN2(n72), .IN3(n128), .Q(n70) );
  AO221X1 U25 ( .IN1(N232), .IN2(n128), .IN3(diff[9]), .IN4(n131), .IN5(n74), 
        .Q(wr_data[9]) );
  AO22X1 U26 ( .IN1(data_in[9]), .IN2(n133), .IN3(N200), .IN4(n135), .Q(n74)
         );
  AO221X1 U27 ( .IN1(N231), .IN2(n128), .IN3(diff[8]), .IN4(n131), .IN5(n75), 
        .Q(wr_data[8]) );
  AO22X1 U28 ( .IN1(data_in[8]), .IN2(n134), .IN3(N199), .IN4(n135), .Q(n75)
         );
  AO221X1 U29 ( .IN1(N230), .IN2(n128), .IN3(diff[7]), .IN4(n131), .IN5(n76), 
        .Q(wr_data[7]) );
  AO22X1 U30 ( .IN1(data_in[7]), .IN2(n134), .IN3(N198), .IN4(n135), .Q(n76)
         );
  AO221X1 U31 ( .IN1(N229), .IN2(n128), .IN3(diff[6]), .IN4(n131), .IN5(n77), 
        .Q(wr_data[6]) );
  AO22X1 U32 ( .IN1(data_in[6]), .IN2(n134), .IN3(N197), .IN4(n135), .Q(n77)
         );
  AO221X1 U33 ( .IN1(N228), .IN2(n128), .IN3(diff[5]), .IN4(n131), .IN5(n78), 
        .Q(wr_data[5]) );
  AO22X1 U34 ( .IN1(data_in[5]), .IN2(n134), .IN3(N196), .IN4(n135), .Q(n78)
         );
  AO221X1 U35 ( .IN1(N227), .IN2(n128), .IN3(diff[4]), .IN4(n131), .IN5(n79), 
        .Q(wr_data[4]) );
  AO22X1 U36 ( .IN1(data_in[4]), .IN2(n134), .IN3(N195), .IN4(n135), .Q(n79)
         );
  AO221X1 U37 ( .IN1(N226), .IN2(n128), .IN3(diff[3]), .IN4(n131), .IN5(n80), 
        .Q(wr_data[3]) );
  AO22X1 U38 ( .IN1(data_in[3]), .IN2(n134), .IN3(N194), .IN4(n135), .Q(n80)
         );
  AO221X1 U39 ( .IN1(N254), .IN2(n128), .IN3(diff[31]), .IN4(n131), .IN5(n81), 
        .Q(wr_data[31]) );
  AO22X1 U40 ( .IN1(data_in[31]), .IN2(n134), .IN3(N222), .IN4(n135), .Q(n81)
         );
  AO221X1 U41 ( .IN1(N253), .IN2(n128), .IN3(diff[30]), .IN4(n131), .IN5(n82), 
        .Q(wr_data[30]) );
  AO22X1 U42 ( .IN1(data_in[30]), .IN2(n134), .IN3(N221), .IN4(n135), .Q(n82)
         );
  AO221X1 U43 ( .IN1(N225), .IN2(n128), .IN3(diff[2]), .IN4(n131), .IN5(n83), 
        .Q(wr_data[2]) );
  AO22X1 U44 ( .IN1(data_in[2]), .IN2(n134), .IN3(N193), .IN4(n135), .Q(n83)
         );
  AO221X1 U45 ( .IN1(N252), .IN2(n128), .IN3(diff[29]), .IN4(n131), .IN5(n84), 
        .Q(wr_data[29]) );
  AO22X1 U46 ( .IN1(data_in[29]), .IN2(n134), .IN3(N220), .IN4(n135), .Q(n84)
         );
  AO221X1 U47 ( .IN1(N251), .IN2(n128), .IN3(diff[28]), .IN4(n131), .IN5(n85), 
        .Q(wr_data[28]) );
  AO22X1 U48 ( .IN1(data_in[28]), .IN2(n134), .IN3(N219), .IN4(n135), .Q(n85)
         );
  AO221X1 U49 ( .IN1(N250), .IN2(n128), .IN3(diff[27]), .IN4(n131), .IN5(n86), 
        .Q(wr_data[27]) );
  AO22X1 U50 ( .IN1(data_in[27]), .IN2(n134), .IN3(N218), .IN4(n135), .Q(n86)
         );
  AO221X1 U51 ( .IN1(N249), .IN2(n129), .IN3(diff[26]), .IN4(n131), .IN5(n87), 
        .Q(wr_data[26]) );
  AO22X1 U52 ( .IN1(data_in[26]), .IN2(n134), .IN3(N217), .IN4(n135), .Q(n87)
         );
  AO221X1 U53 ( .IN1(N248), .IN2(n129), .IN3(diff[25]), .IN4(n131), .IN5(n88), 
        .Q(wr_data[25]) );
  AO22X1 U54 ( .IN1(data_in[25]), .IN2(n134), .IN3(N216), .IN4(n135), .Q(n88)
         );
  AO221X1 U55 ( .IN1(N247), .IN2(n129), .IN3(diff[24]), .IN4(n131), .IN5(n89), 
        .Q(wr_data[24]) );
  AO22X1 U56 ( .IN1(data_in[24]), .IN2(n133), .IN3(N215), .IN4(n135), .Q(n89)
         );
  AO221X1 U57 ( .IN1(N246), .IN2(n129), .IN3(diff[23]), .IN4(n132), .IN5(n90), 
        .Q(wr_data[23]) );
  AO22X1 U58 ( .IN1(data_in[23]), .IN2(n133), .IN3(N214), .IN4(n135), .Q(n90)
         );
  AO221X1 U59 ( .IN1(N245), .IN2(n129), .IN3(diff[22]), .IN4(n132), .IN5(n91), 
        .Q(wr_data[22]) );
  AO22X1 U60 ( .IN1(data_in[22]), .IN2(n133), .IN3(N213), .IN4(n135), .Q(n91)
         );
  AO221X1 U61 ( .IN1(N244), .IN2(n129), .IN3(diff[21]), .IN4(n132), .IN5(n92), 
        .Q(wr_data[21]) );
  AO22X1 U62 ( .IN1(data_in[21]), .IN2(n133), .IN3(N212), .IN4(n136), .Q(n92)
         );
  AO221X1 U63 ( .IN1(N243), .IN2(n129), .IN3(diff[20]), .IN4(n132), .IN5(n93), 
        .Q(wr_data[20]) );
  AO22X1 U64 ( .IN1(data_in[20]), .IN2(n133), .IN3(N211), .IN4(n136), .Q(n93)
         );
  AO221X1 U65 ( .IN1(N224), .IN2(n129), .IN3(diff[1]), .IN4(n132), .IN5(n94), 
        .Q(wr_data[1]) );
  AO22X1 U66 ( .IN1(data_in[1]), .IN2(n133), .IN3(N192), .IN4(n136), .Q(n94)
         );
  AO221X1 U67 ( .IN1(N242), .IN2(n129), .IN3(diff[19]), .IN4(n132), .IN5(n95), 
        .Q(wr_data[19]) );
  AO22X1 U68 ( .IN1(data_in[19]), .IN2(n133), .IN3(N210), .IN4(n136), .Q(n95)
         );
  AO221X1 U69 ( .IN1(N241), .IN2(n129), .IN3(diff[18]), .IN4(n132), .IN5(n96), 
        .Q(wr_data[18]) );
  AO22X1 U70 ( .IN1(data_in[18]), .IN2(n133), .IN3(N209), .IN4(n136), .Q(n96)
         );
  AO221X1 U71 ( .IN1(N240), .IN2(n129), .IN3(diff[17]), .IN4(n132), .IN5(n97), 
        .Q(wr_data[17]) );
  AO22X1 U72 ( .IN1(data_in[17]), .IN2(n133), .IN3(N208), .IN4(n136), .Q(n97)
         );
  AO221X1 U73 ( .IN1(N239), .IN2(n129), .IN3(diff[16]), .IN4(n132), .IN5(n98), 
        .Q(wr_data[16]) );
  AO22X1 U74 ( .IN1(data_in[16]), .IN2(n133), .IN3(N207), .IN4(n136), .Q(n98)
         );
  AO221X1 U75 ( .IN1(N238), .IN2(n129), .IN3(diff[15]), .IN4(n132), .IN5(n99), 
        .Q(wr_data[15]) );
  AO22X1 U76 ( .IN1(data_in[15]), .IN2(n133), .IN3(N206), .IN4(n136), .Q(n99)
         );
  AO221X1 U77 ( .IN1(N237), .IN2(n129), .IN3(diff[14]), .IN4(n132), .IN5(n100), 
        .Q(wr_data[14]) );
  AO22X1 U78 ( .IN1(data_in[14]), .IN2(n133), .IN3(N205), .IN4(n136), .Q(n100)
         );
  AO221X1 U79 ( .IN1(N236), .IN2(n130), .IN3(diff[13]), .IN4(n132), .IN5(n101), 
        .Q(wr_data[13]) );
  AO22X1 U80 ( .IN1(data_in[13]), .IN2(n133), .IN3(N204), .IN4(n136), .Q(n101)
         );
  AO221X1 U81 ( .IN1(N235), .IN2(n130), .IN3(diff[12]), .IN4(n132), .IN5(n102), 
        .Q(wr_data[12]) );
  AO22X1 U82 ( .IN1(data_in[12]), .IN2(n133), .IN3(N203), .IN4(n136), .Q(n102)
         );
  AO221X1 U83 ( .IN1(N234), .IN2(n130), .IN3(diff[11]), .IN4(n132), .IN5(n103), 
        .Q(wr_data[11]) );
  AO22X1 U84 ( .IN1(data_in[11]), .IN2(n133), .IN3(N202), .IN4(n136), .Q(n103)
         );
  AO221X1 U85 ( .IN1(N233), .IN2(n130), .IN3(diff[10]), .IN4(n132), .IN5(n104), 
        .Q(wr_data[10]) );
  AO22X1 U86 ( .IN1(data_in[10]), .IN2(n133), .IN3(N201), .IN4(n136), .Q(n104)
         );
  AO221X1 U87 ( .IN1(N191), .IN2(n136), .IN3(data_in[0]), .IN4(n133), .IN5(
        n105), .Q(wr_data[0]) );
  AO221X1 U88 ( .IN1(N223), .IN2(n130), .IN3(diff[0]), .IN4(n132), .IN5(n106), 
        .Q(n105) );
  AND3X1 U89 ( .IN1(n71), .IN2(n107), .IN3(n72), .Q(n106) );
  AO22X1 U90 ( .IN1(\diff_immed[31] ), .IN2(n158), .IN3(diff[31]), .IN4(
        inst[5]), .Q(n107) );
  AND2X1 U91 ( .IN1(n109), .IN2(n71), .Q(n73) );
  AO22X1 U92 ( .IN1(inst[20]), .IN2(n111), .IN3(n137), .IN4(n112), .Q(
        wr_addr[4]) );
  AO22X1 U93 ( .IN1(inst[19]), .IN2(n111), .IN3(inst[14]), .IN4(n112), .Q(
        wr_addr[3]) );
  AO22X1 U94 ( .IN1(inst[18]), .IN2(n111), .IN3(inst[13]), .IN4(n112), .Q(
        wr_addr[2]) );
  AO22X1 U95 ( .IN1(inst[17]), .IN2(n111), .IN3(inst[12]), .IN4(n112), .Q(
        wr_addr[1]) );
  AO22X1 U96 ( .IN1(inst[16]), .IN2(n111), .IN3(inst[11]), .IN4(n112), .Q(
        wr_addr[0]) );
  AND2X1 U97 ( .IN1(n71), .IN2(n113), .Q(n112) );
  NAND3X0 U98 ( .IN1(n108), .IN2(n110), .IN3(n114), .QN(n113) );
  NAND3X0 U99 ( .IN1(n160), .IN2(n159), .IN3(inst[5]), .QN(n110) );
  NAND3X0 U100 ( .IN1(inst[5]), .IN2(n159), .IN3(inst[1]), .QN(n108) );
  AO21X1 U101 ( .IN1(n71), .IN2(n115), .IN3(n133), .Q(n111) );
  AO21X1 U102 ( .IN1(n72), .IN2(n158), .IN3(n109), .Q(n115) );
  NOR3X0 U103 ( .IN1(inst[1]), .IN2(inst[5]), .IN3(n159), .QN(n109) );
  NOR4X0 U104 ( .IN1(inst[26]), .IN2(inst[0]), .IN3(n117), .IN4(n118), .QN(n71) );
  OR4X1 U105 ( .IN1(inst[2]), .IN2(inst[27]), .IN3(inst[4]), .IN4(inst[31]), 
        .Q(n118) );
  OR3X1 U106 ( .IN1(inst[29]), .IN2(inst[30]), .IN3(inst[28]), .Q(n117) );
  NOR4X0 U107 ( .IN1(inst[30]), .IN2(inst[28]), .IN3(n116), .IN4(n156), .QN(
        data_wr) );
  NAND3X0 U108 ( .IN1(inst[27]), .IN2(inst[26]), .IN3(inst[31]), .QN(n116) );
  AO22X1 U109 ( .IN1(N86), .IN2(n125), .IN3(N54), .IN4(n119), .Q(N150) );
  AO22X1 U110 ( .IN1(N85), .IN2(n125), .IN3(N53), .IN4(n119), .Q(N149) );
  AO22X1 U111 ( .IN1(N84), .IN2(n125), .IN3(N52), .IN4(n119), .Q(N148) );
  AO22X1 U112 ( .IN1(N83), .IN2(n125), .IN3(N51), .IN4(n119), .Q(N147) );
  AO22X1 U113 ( .IN1(N82), .IN2(n126), .IN3(N50), .IN4(n119), .Q(N146) );
  AO22X1 U114 ( .IN1(N81), .IN2(n127), .IN3(N49), .IN4(n119), .Q(N145) );
  AO22X1 U115 ( .IN1(N80), .IN2(n127), .IN3(N48), .IN4(n119), .Q(N144) );
  AO22X1 U116 ( .IN1(N79), .IN2(n126), .IN3(N47), .IN4(n119), .Q(N143) );
  AO22X1 U117 ( .IN1(N78), .IN2(n127), .IN3(N46), .IN4(n124), .Q(N142) );
  AO22X1 U118 ( .IN1(N77), .IN2(n127), .IN3(N45), .IN4(n124), .Q(N141) );
  AO22X1 U119 ( .IN1(N76), .IN2(n126), .IN3(N44), .IN4(n124), .Q(N140) );
  AO22X1 U120 ( .IN1(N75), .IN2(n126), .IN3(N43), .IN4(n124), .Q(N139) );
  AO22X1 U121 ( .IN1(N74), .IN2(n126), .IN3(N42), .IN4(n124), .Q(N138) );
  AO22X1 U122 ( .IN1(N73), .IN2(n126), .IN3(N41), .IN4(n124), .Q(N137) );
  AO22X1 U123 ( .IN1(N72), .IN2(n126), .IN3(N40), .IN4(n124), .Q(N136) );
  AO22X1 U124 ( .IN1(N71), .IN2(n126), .IN3(N39), .IN4(n124), .Q(N135) );
  AO22X1 U125 ( .IN1(N70), .IN2(n126), .IN3(N38), .IN4(n124), .Q(N134) );
  AO22X1 U126 ( .IN1(N69), .IN2(n126), .IN3(N37), .IN4(n124), .Q(N133) );
  AO22X1 U127 ( .IN1(N68), .IN2(n126), .IN3(N36), .IN4(n124), .Q(N132) );
  AO22X1 U128 ( .IN1(N67), .IN2(n127), .IN3(N35), .IN4(n124), .Q(N131) );
  AO22X1 U129 ( .IN1(N66), .IN2(n126), .IN3(N34), .IN4(n123), .Q(N130) );
  AO22X1 U130 ( .IN1(N65), .IN2(n127), .IN3(N33), .IN4(n123), .Q(N129) );
  AO22X1 U131 ( .IN1(N64), .IN2(n126), .IN3(N32), .IN4(n123), .Q(N128) );
  AO22X1 U132 ( .IN1(N63), .IN2(n127), .IN3(N31), .IN4(n123), .Q(N127) );
  AO22X1 U133 ( .IN1(N62), .IN2(n126), .IN3(N30), .IN4(n123), .Q(N126) );
  AO22X1 U134 ( .IN1(N61), .IN2(n127), .IN3(N29), .IN4(n123), .Q(N125) );
  AO22X1 U135 ( .IN1(N60), .IN2(n127), .IN3(N28), .IN4(n123), .Q(N124) );
  AO22X1 U136 ( .IN1(N59), .IN2(n127), .IN3(N27), .IN4(n123), .Q(N123) );
  AO22X1 U137 ( .IN1(N58), .IN2(n127), .IN3(N26), .IN4(n123), .Q(N122) );
  AO22X1 U138 ( .IN1(N57), .IN2(n127), .IN3(N25), .IN4(n123), .Q(N121) );
  AO22X1 U139 ( .IN1(N56), .IN2(n127), .IN3(N24), .IN4(n123), .Q(N120) );
  AO22X1 U140 ( .IN1(N55), .IN2(n127), .IN3(N23), .IN4(n123), .Q(N119) );
  NAND4X0 U141 ( .IN1(N378), .IN2(n157), .IN3(inst[28]), .IN4(n120), .QN(n119)
         );
  NOR3X0 U142 ( .IN1(inst[29]), .IN2(inst[31]), .IN3(inst[30]), .QN(n120) );
  regfile RF ( .clk(clk), .nrst(n143), .rd_addrA(inst[25:21]), .rd_addrB(
        inst[20:16]), .wr_addr(wr_addr), .wr_en(wr_en), .wr_data(wr_data), 
        .rd_dataA(rd_dataA), .rd_dataB(data_out) );
  single_cycle_mips_DW01_add_0 add_123 ( .A(rd_dataA), .B({n139, n139, n138, 
        n139, n139, n139, n139, n138, n138, n138, n138, n138, n137, n137, n137, 
        n137, n137, inst[14:0]}), .CI(1'b0), .SUM(data_addr) );
  single_cycle_mips_DW01_add_1 add_91 ( .A(rd_dataA), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n137, inst[14:0]}), .CI(1'b0), .SUM({N254, N253, N252, N251, 
        N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, 
        N238, N237, N236, N235, N234, N233, N232, N231, N230, N229, N228, N227, 
        N226, N225, N224, N223}) );
  single_cycle_mips_DW01_add_2 add_70 ( .A(rd_dataA), .B(data_out), .CI(1'b0), 
        .SUM({N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202, N201, N200, 
        N199, N198, N197, N196, N195, N194, N193, N192, N191}) );
  single_cycle_mips_DW01_sub_0 sub_63 ( .A(rd_dataA), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, n138, inst[14:0]}), .CI(1'b0), .DIFF({\diff_immed[31] , 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30}) );
  single_cycle_mips_DW01_add_3 add_0_root_add_25_2 ( .A({n140, n140, n140, 
        n140, n140, n140, n141, n141, n141, n141, n141, n141, n141, n142, n142, 
        n142, n140, inst[14:0]}), .B({N54, N53, N52, N51, N50, N49, N48, N47, 
        N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, 
        N32, N31, N30, N29, N28, N27, N26, N25, N24, N23}), .CI(1'b0), .SUM({
        N86, N85, N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, 
        N72, N71, N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, 
        N58, N57, N56, N55}) );
  single_cycle_mips_DW01_add_4 r102 ( .A(inst_addr), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N54, N53, N52, N51, 
        N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, 
        N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, N26, N25, N24, N23})
         );
  single_cycle_mips_DW01_sub_1 sub_62 ( .A(rd_dataA), .B({data_out[15], 
        data_out[15], data_out[15], data_out[15], data_out[15], data_out[15], 
        data_out[15], data_out[15], data_out[15], data_out[15], data_out[15], 
        data_out[15], data_out[15], data_out[15], data_out[15], data_out[15], 
        data_out[15:0]}), .CI(1'b0), .DIFF(diff) );
  NBUFFX2 U143 ( .INP(n67), .Z(n135) );
  NBUFFX2 U144 ( .INP(n69), .Z(n131) );
  NBUFFX2 U145 ( .INP(n68), .Z(n133) );
  NBUFFX2 U146 ( .INP(n73), .Z(n128) );
  NBUFFX2 U147 ( .INP(n69), .Z(n132) );
  NBUFFX2 U148 ( .INP(n67), .Z(n136) );
  NBUFFX2 U149 ( .INP(n73), .Z(n129) );
  NBUFFX2 U150 ( .INP(n68), .Z(n134) );
  NBUFFX2 U151 ( .INP(n73), .Z(n130) );
  INVX0 U152 ( .INP(n119), .ZN(n125) );
  INVX0 U153 ( .INP(n119), .ZN(n126) );
  INVX0 U154 ( .INP(n119), .ZN(n127) );
  INVX0 U155 ( .INP(n71), .ZN(n155) );
  NOR2X0 U156 ( .IN1(n155), .IN2(n110), .QN(n67) );
  NOR2X0 U157 ( .IN1(n108), .IN2(n155), .QN(n69) );
  NOR2X0 U158 ( .IN1(n159), .IN2(n160), .QN(n72) );
  NOR2X0 U159 ( .IN1(n116), .IN2(n117), .QN(n68) );
  NBUFFX4 U160 ( .INP(n143), .Z(n122) );
  INVX0 U161 ( .INP(inst[27]), .ZN(n157) );
  NBUFFX4 U162 ( .INP(inst[15]), .Z(n137) );
  NBUFFX4 U163 ( .INP(inst[15]), .Z(n138) );
  NBUFFX4 U164 ( .INP(inst[15]), .Z(n139) );
  INVX0 U165 ( .INP(inst[29]), .ZN(n156) );
  INVX0 U166 ( .INP(inst[3]), .ZN(n159) );
  INVX0 U167 ( .INP(inst[1]), .ZN(n160) );
  NAND2X1 U168 ( .IN1(n72), .IN2(inst[5]), .QN(n114) );
  INVX0 U169 ( .INP(inst[5]), .ZN(n158) );
  NBUFFX4 U170 ( .INP(inst[15]), .Z(n140) );
  NBUFFX4 U171 ( .INP(inst[15]), .Z(n141) );
  NBUFFX2 U172 ( .INP(inst[15]), .Z(n142) );
  NBUFFX4 U173 ( .INP(rst_n), .Z(n144) );
  NBUFFX2 U174 ( .INP(rst_n), .Z(n143) );
  INVX0 U175 ( .INP(n125), .ZN(n123) );
  INVX0 U176 ( .INP(n125), .ZN(n124) );
  NOR4X0 U177 ( .IN1(diff[27]), .IN2(diff[26]), .IN3(diff[25]), .IN4(diff[24]), 
        .QN(n148) );
  NOR4X0 U178 ( .IN1(diff[30]), .IN2(diff[2]), .IN3(diff[29]), .IN4(diff[28]), 
        .QN(n147) );
  NOR4X0 U179 ( .IN1(diff[5]), .IN2(diff[4]), .IN3(diff[3]), .IN4(diff[31]), 
        .QN(n146) );
  NOR4X0 U180 ( .IN1(diff[9]), .IN2(diff[8]), .IN3(diff[7]), .IN4(diff[6]), 
        .QN(n145) );
  NAND4X0 U181 ( .IN1(n148), .IN2(n147), .IN3(n146), .IN4(n145), .QN(n154) );
  NOR4X0 U182 ( .IN1(diff[12]), .IN2(diff[11]), .IN3(diff[10]), .IN4(diff[0]), 
        .QN(n152) );
  NOR4X0 U183 ( .IN1(diff[16]), .IN2(diff[15]), .IN3(diff[14]), .IN4(diff[13]), 
        .QN(n151) );
  NOR4X0 U184 ( .IN1(diff[1]), .IN2(diff[19]), .IN3(diff[18]), .IN4(diff[17]), 
        .QN(n150) );
  NOR4X0 U185 ( .IN1(diff[23]), .IN2(diff[22]), .IN3(diff[21]), .IN4(diff[20]), 
        .QN(n149) );
  NAND4X0 U186 ( .IN1(n152), .IN2(n151), .IN3(n150), .IN4(n149), .QN(n153) );
  NOR2X0 U187 ( .IN1(n154), .IN2(n153), .QN(N378) );
endmodule

