`timescale 1ns/1ps
module rf ( clk, nrst, rd_addrA, rd_addrB, rd_dataA, rd_dataB, wr_en, wr_addr, 
        wr_data );
  input [4:0] rd_addrA;
  input [4:0] rd_addrB;
  output [31:0] rd_dataA;
  output [31:0] rd_dataB;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  input clk, nrst, wr_en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, \regf[31][31] ,
         \regf[31][30] , \regf[31][29] , \regf[31][28] , \regf[31][27] ,
         \regf[31][26] , \regf[31][25] , \regf[31][24] , \regf[31][23] ,
         \regf[31][22] , \regf[31][21] , \regf[31][20] , \regf[31][19] ,
         \regf[31][18] , \regf[31][17] , \regf[31][16] , \regf[31][15] ,
         \regf[31][14] , \regf[31][13] , \regf[31][12] , \regf[31][11] ,
         \regf[31][10] , \regf[31][9] , \regf[31][8] , \regf[31][7] ,
         \regf[31][6] , \regf[31][5] , \regf[31][4] , \regf[31][3] ,
         \regf[31][2] , \regf[31][1] , \regf[31][0] , \regf[30][31] ,
         \regf[30][30] , \regf[30][29] , \regf[30][28] , \regf[30][27] ,
         \regf[30][26] , \regf[30][25] , \regf[30][24] , \regf[30][23] ,
         \regf[30][22] , \regf[30][21] , \regf[30][20] , \regf[30][19] ,
         \regf[30][18] , \regf[30][17] , \regf[30][16] , \regf[30][15] ,
         \regf[30][14] , \regf[30][13] , \regf[30][12] , \regf[30][11] ,
         \regf[30][10] , \regf[30][9] , \regf[30][8] , \regf[30][7] ,
         \regf[30][6] , \regf[30][5] , \regf[30][4] , \regf[30][3] ,
         \regf[30][2] , \regf[30][1] , \regf[30][0] , \regf[29][31] ,
         \regf[29][30] , \regf[29][29] , \regf[29][28] , \regf[29][27] ,
         \regf[29][26] , \regf[29][25] , \regf[29][24] , \regf[29][23] ,
         \regf[29][22] , \regf[29][21] , \regf[29][20] , \regf[29][19] ,
         \regf[29][18] , \regf[29][17] , \regf[29][16] , \regf[29][15] ,
         \regf[29][14] , \regf[29][13] , \regf[29][12] , \regf[29][11] ,
         \regf[29][10] , \regf[29][9] , \regf[29][8] , \regf[29][7] ,
         \regf[29][6] , \regf[29][5] , \regf[29][4] , \regf[29][3] ,
         \regf[29][2] , \regf[29][1] , \regf[29][0] , \regf[28][31] ,
         \regf[28][30] , \regf[28][29] , \regf[28][28] , \regf[28][27] ,
         \regf[28][26] , \regf[28][25] , \regf[28][24] , \regf[28][23] ,
         \regf[28][22] , \regf[28][21] , \regf[28][20] , \regf[28][19] ,
         \regf[28][18] , \regf[28][17] , \regf[28][16] , \regf[28][15] ,
         \regf[28][14] , \regf[28][13] , \regf[28][12] , \regf[28][11] ,
         \regf[28][10] , \regf[28][9] , \regf[28][8] , \regf[28][7] ,
         \regf[28][6] , \regf[28][5] , \regf[28][4] , \regf[28][3] ,
         \regf[28][2] , \regf[28][1] , \regf[28][0] , \regf[27][31] ,
         \regf[27][30] , \regf[27][29] , \regf[27][28] , \regf[27][27] ,
         \regf[27][26] , \regf[27][25] , \regf[27][24] , \regf[27][23] ,
         \regf[27][22] , \regf[27][21] , \regf[27][20] , \regf[27][19] ,
         \regf[27][18] , \regf[27][17] , \regf[27][16] , \regf[27][15] ,
         \regf[27][14] , \regf[27][13] , \regf[27][12] , \regf[27][11] ,
         \regf[27][10] , \regf[27][9] , \regf[27][8] , \regf[27][7] ,
         \regf[27][6] , \regf[27][5] , \regf[27][4] , \regf[27][3] ,
         \regf[27][2] , \regf[27][1] , \regf[27][0] , \regf[26][31] ,
         \regf[26][30] , \regf[26][29] , \regf[26][28] , \regf[26][27] ,
         \regf[26][26] , \regf[26][25] , \regf[26][24] , \regf[26][23] ,
         \regf[26][22] , \regf[26][21] , \regf[26][20] , \regf[26][19] ,
         \regf[26][18] , \regf[26][17] , \regf[26][16] , \regf[26][15] ,
         \regf[26][14] , \regf[26][13] , \regf[26][12] , \regf[26][11] ,
         \regf[26][10] , \regf[26][9] , \regf[26][8] , \regf[26][7] ,
         \regf[26][6] , \regf[26][5] , \regf[26][4] , \regf[26][3] ,
         \regf[26][2] , \regf[26][1] , \regf[26][0] , \regf[25][31] ,
         \regf[25][30] , \regf[25][29] , \regf[25][28] , \regf[25][27] ,
         \regf[25][26] , \regf[25][25] , \regf[25][24] , \regf[25][23] ,
         \regf[25][22] , \regf[25][21] , \regf[25][20] , \regf[25][19] ,
         \regf[25][18] , \regf[25][17] , \regf[25][16] , \regf[25][15] ,
         \regf[25][14] , \regf[25][13] , \regf[25][12] , \regf[25][11] ,
         \regf[25][10] , \regf[25][9] , \regf[25][8] , \regf[25][7] ,
         \regf[25][6] , \regf[25][5] , \regf[25][4] , \regf[25][3] ,
         \regf[25][2] , \regf[25][1] , \regf[25][0] , \regf[24][31] ,
         \regf[24][30] , \regf[24][29] , \regf[24][28] , \regf[24][27] ,
         \regf[24][26] , \regf[24][25] , \regf[24][24] , \regf[24][23] ,
         \regf[24][22] , \regf[24][21] , \regf[24][20] , \regf[24][19] ,
         \regf[24][18] , \regf[24][17] , \regf[24][16] , \regf[24][15] ,
         \regf[24][14] , \regf[24][13] , \regf[24][12] , \regf[24][11] ,
         \regf[24][10] , \regf[24][9] , \regf[24][8] , \regf[24][7] ,
         \regf[24][6] , \regf[24][5] , \regf[24][4] , \regf[24][3] ,
         \regf[24][2] , \regf[24][1] , \regf[24][0] , \regf[23][31] ,
         \regf[23][30] , \regf[23][29] , \regf[23][28] , \regf[23][27] ,
         \regf[23][26] , \regf[23][25] , \regf[23][24] , \regf[23][23] ,
         \regf[23][22] , \regf[23][21] , \regf[23][20] , \regf[23][19] ,
         \regf[23][18] , \regf[23][17] , \regf[23][16] , \regf[23][15] ,
         \regf[23][14] , \regf[23][13] , \regf[23][12] , \regf[23][11] ,
         \regf[23][10] , \regf[23][9] , \regf[23][8] , \regf[23][7] ,
         \regf[23][6] , \regf[23][5] , \regf[23][4] , \regf[23][3] ,
         \regf[23][2] , \regf[23][1] , \regf[23][0] , \regf[22][31] ,
         \regf[22][30] , \regf[22][29] , \regf[22][28] , \regf[22][27] ,
         \regf[22][26] , \regf[22][25] , \regf[22][24] , \regf[22][23] ,
         \regf[22][22] , \regf[22][21] , \regf[22][20] , \regf[22][19] ,
         \regf[22][18] , \regf[22][17] , \regf[22][16] , \regf[22][15] ,
         \regf[22][14] , \regf[22][13] , \regf[22][12] , \regf[22][11] ,
         \regf[22][10] , \regf[22][9] , \regf[22][8] , \regf[22][7] ,
         \regf[22][6] , \regf[22][5] , \regf[22][4] , \regf[22][3] ,
         \regf[22][2] , \regf[22][1] , \regf[22][0] , \regf[21][31] ,
         \regf[21][30] , \regf[21][29] , \regf[21][28] , \regf[21][27] ,
         \regf[21][26] , \regf[21][25] , \regf[21][24] , \regf[21][23] ,
         \regf[21][22] , \regf[21][21] , \regf[21][20] , \regf[21][19] ,
         \regf[21][18] , \regf[21][17] , \regf[21][16] , \regf[21][15] ,
         \regf[21][14] , \regf[21][13] , \regf[21][12] , \regf[21][11] ,
         \regf[21][10] , \regf[21][9] , \regf[21][8] , \regf[21][7] ,
         \regf[21][6] , \regf[21][5] , \regf[21][4] , \regf[21][3] ,
         \regf[21][2] , \regf[21][1] , \regf[21][0] , \regf[20][31] ,
         \regf[20][30] , \regf[20][29] , \regf[20][28] , \regf[20][27] ,
         \regf[20][26] , \regf[20][25] , \regf[20][24] , \regf[20][23] ,
         \regf[20][22] , \regf[20][21] , \regf[20][20] , \regf[20][19] ,
         \regf[20][18] , \regf[20][17] , \regf[20][16] , \regf[20][15] ,
         \regf[20][14] , \regf[20][13] , \regf[20][12] , \regf[20][11] ,
         \regf[20][10] , \regf[20][9] , \regf[20][8] , \regf[20][7] ,
         \regf[20][6] , \regf[20][5] , \regf[20][4] , \regf[20][3] ,
         \regf[20][2] , \regf[20][1] , \regf[20][0] , \regf[19][31] ,
         \regf[19][30] , \regf[19][29] , \regf[19][28] , \regf[19][27] ,
         \regf[19][26] , \regf[19][25] , \regf[19][24] , \regf[19][23] ,
         \regf[19][22] , \regf[19][21] , \regf[19][20] , \regf[19][19] ,
         \regf[19][18] , \regf[19][17] , \regf[19][16] , \regf[19][15] ,
         \regf[19][14] , \regf[19][13] , \regf[19][12] , \regf[19][11] ,
         \regf[19][10] , \regf[19][9] , \regf[19][8] , \regf[19][7] ,
         \regf[19][6] , \regf[19][5] , \regf[19][4] , \regf[19][3] ,
         \regf[19][2] , \regf[19][1] , \regf[19][0] , \regf[18][31] ,
         \regf[18][30] , \regf[18][29] , \regf[18][28] , \regf[18][27] ,
         \regf[18][26] , \regf[18][25] , \regf[18][24] , \regf[18][23] ,
         \regf[18][22] , \regf[18][21] , \regf[18][20] , \regf[18][19] ,
         \regf[18][18] , \regf[18][17] , \regf[18][16] , \regf[18][15] ,
         \regf[18][14] , \regf[18][13] , \regf[18][12] , \regf[18][11] ,
         \regf[18][10] , \regf[18][9] , \regf[18][8] , \regf[18][7] ,
         \regf[18][6] , \regf[18][5] , \regf[18][4] , \regf[18][3] ,
         \regf[18][2] , \regf[18][1] , \regf[18][0] , \regf[17][31] ,
         \regf[17][30] , \regf[17][29] , \regf[17][28] , \regf[17][27] ,
         \regf[17][26] , \regf[17][25] , \regf[17][24] , \regf[17][23] ,
         \regf[17][22] , \regf[17][21] , \regf[17][20] , \regf[17][19] ,
         \regf[17][18] , \regf[17][17] , \regf[17][16] , \regf[17][15] ,
         \regf[17][14] , \regf[17][13] , \regf[17][12] , \regf[17][11] ,
         \regf[17][10] , \regf[17][9] , \regf[17][8] , \regf[17][7] ,
         \regf[17][6] , \regf[17][5] , \regf[17][4] , \regf[17][3] ,
         \regf[17][2] , \regf[17][1] , \regf[17][0] , \regf[16][31] ,
         \regf[16][30] , \regf[16][29] , \regf[16][28] , \regf[16][27] ,
         \regf[16][26] , \regf[16][25] , \regf[16][24] , \regf[16][23] ,
         \regf[16][22] , \regf[16][21] , \regf[16][20] , \regf[16][19] ,
         \regf[16][18] , \regf[16][17] , \regf[16][16] , \regf[16][15] ,
         \regf[16][14] , \regf[16][13] , \regf[16][12] , \regf[16][11] ,
         \regf[16][10] , \regf[16][9] , \regf[16][8] , \regf[16][7] ,
         \regf[16][6] , \regf[16][5] , \regf[16][4] , \regf[16][3] ,
         \regf[16][2] , \regf[16][1] , \regf[16][0] , \regf[15][31] ,
         \regf[15][30] , \regf[15][29] , \regf[15][28] , \regf[15][27] ,
         \regf[15][26] , \regf[15][25] , \regf[15][24] , \regf[15][23] ,
         \regf[15][22] , \regf[15][21] , \regf[15][20] , \regf[15][19] ,
         \regf[15][18] , \regf[15][17] , \regf[15][16] , \regf[15][15] ,
         \regf[15][14] , \regf[15][13] , \regf[15][12] , \regf[15][11] ,
         \regf[15][10] , \regf[15][9] , \regf[15][8] , \regf[15][7] ,
         \regf[15][6] , \regf[15][5] , \regf[15][4] , \regf[15][3] ,
         \regf[15][2] , \regf[15][1] , \regf[15][0] , \regf[14][31] ,
         \regf[14][30] , \regf[14][29] , \regf[14][28] , \regf[14][27] ,
         \regf[14][26] , \regf[14][25] , \regf[14][24] , \regf[14][23] ,
         \regf[14][22] , \regf[14][21] , \regf[14][20] , \regf[14][19] ,
         \regf[14][18] , \regf[14][17] , \regf[14][16] , \regf[14][15] ,
         \regf[14][14] , \regf[14][13] , \regf[14][12] , \regf[14][11] ,
         \regf[14][10] , \regf[14][9] , \regf[14][8] , \regf[14][7] ,
         \regf[14][6] , \regf[14][5] , \regf[14][4] , \regf[14][3] ,
         \regf[14][2] , \regf[14][1] , \regf[14][0] , \regf[13][31] ,
         \regf[13][30] , \regf[13][29] , \regf[13][28] , \regf[13][27] ,
         \regf[13][26] , \regf[13][25] , \regf[13][24] , \regf[13][23] ,
         \regf[13][22] , \regf[13][21] , \regf[13][20] , \regf[13][19] ,
         \regf[13][18] , \regf[13][17] , \regf[13][16] , \regf[13][15] ,
         \regf[13][14] , \regf[13][13] , \regf[13][12] , \regf[13][11] ,
         \regf[13][10] , \regf[13][9] , \regf[13][8] , \regf[13][7] ,
         \regf[13][6] , \regf[13][5] , \regf[13][4] , \regf[13][3] ,
         \regf[13][2] , \regf[13][1] , \regf[13][0] , \regf[12][31] ,
         \regf[12][30] , \regf[12][29] , \regf[12][28] , \regf[12][27] ,
         \regf[12][26] , \regf[12][25] , \regf[12][24] , \regf[12][23] ,
         \regf[12][22] , \regf[12][21] , \regf[12][20] , \regf[12][19] ,
         \regf[12][18] , \regf[12][17] , \regf[12][16] , \regf[12][15] ,
         \regf[12][14] , \regf[12][13] , \regf[12][12] , \regf[12][11] ,
         \regf[12][10] , \regf[12][9] , \regf[12][8] , \regf[12][7] ,
         \regf[12][6] , \regf[12][5] , \regf[12][4] , \regf[12][3] ,
         \regf[12][2] , \regf[12][1] , \regf[12][0] , \regf[11][31] ,
         \regf[11][30] , \regf[11][29] , \regf[11][28] , \regf[11][27] ,
         \regf[11][26] , \regf[11][25] , \regf[11][24] , \regf[11][23] ,
         \regf[11][22] , \regf[11][21] , \regf[11][20] , \regf[11][19] ,
         \regf[11][18] , \regf[11][17] , \regf[11][16] , \regf[11][15] ,
         \regf[11][14] , \regf[11][13] , \regf[11][12] , \regf[11][11] ,
         \regf[11][10] , \regf[11][9] , \regf[11][8] , \regf[11][7] ,
         \regf[11][6] , \regf[11][5] , \regf[11][4] , \regf[11][3] ,
         \regf[11][2] , \regf[11][1] , \regf[11][0] , \regf[10][31] ,
         \regf[10][30] , \regf[10][29] , \regf[10][28] , \regf[10][27] ,
         \regf[10][26] , \regf[10][25] , \regf[10][24] , \regf[10][23] ,
         \regf[10][22] , \regf[10][21] , \regf[10][20] , \regf[10][19] ,
         \regf[10][18] , \regf[10][17] , \regf[10][16] , \regf[10][15] ,
         \regf[10][14] , \regf[10][13] , \regf[10][12] , \regf[10][11] ,
         \regf[10][10] , \regf[10][9] , \regf[10][8] , \regf[10][7] ,
         \regf[10][6] , \regf[10][5] , \regf[10][4] , \regf[10][3] ,
         \regf[10][2] , \regf[10][1] , \regf[10][0] , \regf[9][31] ,
         \regf[9][30] , \regf[9][29] , \regf[9][28] , \regf[9][27] ,
         \regf[9][26] , \regf[9][25] , \regf[9][24] , \regf[9][23] ,
         \regf[9][22] , \regf[9][21] , \regf[9][20] , \regf[9][19] ,
         \regf[9][18] , \regf[9][17] , \regf[9][16] , \regf[9][15] ,
         \regf[9][14] , \regf[9][13] , \regf[9][12] , \regf[9][11] ,
         \regf[9][10] , \regf[9][9] , \regf[9][8] , \regf[9][7] , \regf[9][6] ,
         \regf[9][5] , \regf[9][4] , \regf[9][3] , \regf[9][2] , \regf[9][1] ,
         \regf[9][0] , \regf[8][31] , \regf[8][30] , \regf[8][29] ,
         \regf[8][28] , \regf[8][27] , \regf[8][26] , \regf[8][25] ,
         \regf[8][24] , \regf[8][23] , \regf[8][22] , \regf[8][21] ,
         \regf[8][20] , \regf[8][19] , \regf[8][18] , \regf[8][17] ,
         \regf[8][16] , \regf[8][15] , \regf[8][14] , \regf[8][13] ,
         \regf[8][12] , \regf[8][11] , \regf[8][10] , \regf[8][9] ,
         \regf[8][8] , \regf[8][7] , \regf[8][6] , \regf[8][5] , \regf[8][4] ,
         \regf[8][3] , \regf[8][2] , \regf[8][1] , \regf[8][0] , \regf[7][31] ,
         \regf[7][30] , \regf[7][29] , \regf[7][28] , \regf[7][27] ,
         \regf[7][26] , \regf[7][25] , \regf[7][24] , \regf[7][23] ,
         \regf[7][22] , \regf[7][21] , \regf[7][20] , \regf[7][19] ,
         \regf[7][18] , \regf[7][17] , \regf[7][16] , \regf[7][15] ,
         \regf[7][14] , \regf[7][13] , \regf[7][12] , \regf[7][11] ,
         \regf[7][10] , \regf[7][9] , \regf[7][8] , \regf[7][7] , \regf[7][6] ,
         \regf[7][5] , \regf[7][4] , \regf[7][3] , \regf[7][2] , \regf[7][1] ,
         \regf[7][0] , \regf[6][31] , \regf[6][30] , \regf[6][29] ,
         \regf[6][28] , \regf[6][27] , \regf[6][26] , \regf[6][25] ,
         \regf[6][24] , \regf[6][23] , \regf[6][22] , \regf[6][21] ,
         \regf[6][20] , \regf[6][19] , \regf[6][18] , \regf[6][17] ,
         \regf[6][16] , \regf[6][15] , \regf[6][14] , \regf[6][13] ,
         \regf[6][12] , \regf[6][11] , \regf[6][10] , \regf[6][9] ,
         \regf[6][8] , \regf[6][7] , \regf[6][6] , \regf[6][5] , \regf[6][4] ,
         \regf[6][3] , \regf[6][2] , \regf[6][1] , \regf[6][0] , \regf[5][31] ,
         \regf[5][30] , \regf[5][29] , \regf[5][28] , \regf[5][27] ,
         \regf[5][26] , \regf[5][25] , \regf[5][24] , \regf[5][23] ,
         \regf[5][22] , \regf[5][21] , \regf[5][20] , \regf[5][19] ,
         \regf[5][18] , \regf[5][17] , \regf[5][16] , \regf[5][15] ,
         \regf[5][14] , \regf[5][13] , \regf[5][12] , \regf[5][11] ,
         \regf[5][10] , \regf[5][9] , \regf[5][8] , \regf[5][7] , \regf[5][6] ,
         \regf[5][5] , \regf[5][4] , \regf[5][3] , \regf[5][2] , \regf[5][1] ,
         \regf[5][0] , \regf[4][31] , \regf[4][30] , \regf[4][29] ,
         \regf[4][28] , \regf[4][27] , \regf[4][26] , \regf[4][25] ,
         \regf[4][24] , \regf[4][23] , \regf[4][22] , \regf[4][21] ,
         \regf[4][20] , \regf[4][19] , \regf[4][18] , \regf[4][17] ,
         \regf[4][16] , \regf[4][15] , \regf[4][14] , \regf[4][13] ,
         \regf[4][12] , \regf[4][11] , \regf[4][10] , \regf[4][9] ,
         \regf[4][8] , \regf[4][7] , \regf[4][6] , \regf[4][5] , \regf[4][4] ,
         \regf[4][3] , \regf[4][2] , \regf[4][1] , \regf[4][0] , \regf[3][31] ,
         \regf[3][30] , \regf[3][29] , \regf[3][28] , \regf[3][27] ,
         \regf[3][26] , \regf[3][25] , \regf[3][24] , \regf[3][23] ,
         \regf[3][22] , \regf[3][21] , \regf[3][20] , \regf[3][19] ,
         \regf[3][18] , \regf[3][17] , \regf[3][16] , \regf[3][15] ,
         \regf[3][14] , \regf[3][13] , \regf[3][12] , \regf[3][11] ,
         \regf[3][10] , \regf[3][9] , \regf[3][8] , \regf[3][7] , \regf[3][6] ,
         \regf[3][5] , \regf[3][4] , \regf[3][3] , \regf[3][2] , \regf[3][1] ,
         \regf[3][0] , \regf[2][31] , \regf[2][30] , \regf[2][29] ,
         \regf[2][28] , \regf[2][27] , \regf[2][26] , \regf[2][25] ,
         \regf[2][24] , \regf[2][23] , \regf[2][22] , \regf[2][21] ,
         \regf[2][20] , \regf[2][19] , \regf[2][18] , \regf[2][17] ,
         \regf[2][16] , \regf[2][15] , \regf[2][14] , \regf[2][13] ,
         \regf[2][12] , \regf[2][11] , \regf[2][10] , \regf[2][9] ,
         \regf[2][8] , \regf[2][7] , \regf[2][6] , \regf[2][5] , \regf[2][4] ,
         \regf[2][3] , \regf[2][2] , \regf[2][1] , \regf[2][0] , \regf[1][31] ,
         \regf[1][30] , \regf[1][29] , \regf[1][28] , \regf[1][27] ,
         \regf[1][26] , \regf[1][25] , \regf[1][24] , \regf[1][23] ,
         \regf[1][22] , \regf[1][21] , \regf[1][20] , \regf[1][19] ,
         \regf[1][18] , \regf[1][17] , \regf[1][16] , \regf[1][15] ,
         \regf[1][14] , \regf[1][13] , \regf[1][12] , \regf[1][11] ,
         \regf[1][10] , \regf[1][9] , \regf[1][8] , \regf[1][7] , \regf[1][6] ,
         \regf[1][5] , \regf[1][4] , \regf[1][3] , \regf[1][2] , \regf[1][1] ,
         \regf[1][0] , n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714;
  assign N11 = rd_addrA[0];
  assign N12 = rd_addrA[1];
  assign N13 = rd_addrA[2];
  assign N14 = rd_addrA[3];
  assign N15 = rd_addrA[4];
  assign N16 = rd_addrB[0];
  assign N17 = rd_addrB[1];
  assign N18 = rd_addrB[2];
  assign N19 = rd_addrB[3];
  assign N20 = rd_addrB[4];

  DFFARX1 \regf_reg[31][31]  ( .D(n1070), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][31] ) );
  DFFARX1 \regf_reg[31][30]  ( .D(n1069), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][30] ) );
  DFFARX1 \regf_reg[31][29]  ( .D(n1068), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][29] ) );
  DFFARX1 \regf_reg[31][28]  ( .D(n1067), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][28] ) );
  DFFARX1 \regf_reg[31][27]  ( .D(n1066), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][27] ) );
  DFFARX1 \regf_reg[31][26]  ( .D(n1065), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][26] ) );
  DFFARX1 \regf_reg[31][25]  ( .D(n1064), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][25] ) );
  DFFARX1 \regf_reg[31][24]  ( .D(n1063), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][24] ) );
  DFFARX1 \regf_reg[31][23]  ( .D(n1062), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][23] ) );
  DFFARX1 \regf_reg[31][22]  ( .D(n1061), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][22] ) );
  DFFARX1 \regf_reg[31][21]  ( .D(n1060), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][21] ) );
  DFFARX1 \regf_reg[31][20]  ( .D(n1059), .CLK(clk), .RSTB(n2621), .Q(
        \regf[31][20] ) );
  DFFARX1 \regf_reg[31][19]  ( .D(n1058), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][19] ) );
  DFFARX1 \regf_reg[31][18]  ( .D(n1057), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][18] ) );
  DFFARX1 \regf_reg[31][17]  ( .D(n1056), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][17] ) );
  DFFARX1 \regf_reg[31][16]  ( .D(n1055), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][16] ) );
  DFFARX1 \regf_reg[31][15]  ( .D(n1054), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][15] ) );
  DFFARX1 \regf_reg[31][14]  ( .D(n1053), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][14] ) );
  DFFARX1 \regf_reg[31][13]  ( .D(n1052), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][13] ) );
  DFFARX1 \regf_reg[31][12]  ( .D(n1051), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][12] ) );
  DFFARX1 \regf_reg[31][11]  ( .D(n1050), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][11] ) );
  DFFARX1 \regf_reg[31][10]  ( .D(n1049), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][10] ) );
  DFFARX1 \regf_reg[31][9]  ( .D(n1048), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][9] ) );
  DFFARX1 \regf_reg[31][8]  ( .D(n1047), .CLK(clk), .RSTB(n2622), .Q(
        \regf[31][8] ) );
  DFFARX1 \regf_reg[31][7]  ( .D(n1046), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][7] ) );
  DFFARX1 \regf_reg[31][6]  ( .D(n1045), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][6] ) );
  DFFARX1 \regf_reg[31][5]  ( .D(n1044), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][5] ) );
  DFFARX1 \regf_reg[31][4]  ( .D(n1043), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][4] ) );
  DFFARX1 \regf_reg[31][3]  ( .D(n1042), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][3] ) );
  DFFARX1 \regf_reg[31][2]  ( .D(n1041), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][2] ) );
  DFFARX1 \regf_reg[31][1]  ( .D(n1040), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][1] ) );
  DFFARX1 \regf_reg[31][0]  ( .D(n1039), .CLK(clk), .RSTB(n2623), .Q(
        \regf[31][0] ) );
  DFFARX1 \regf_reg[30][31]  ( .D(n1038), .CLK(clk), .RSTB(n2623), .Q(
        \regf[30][31] ) );
  DFFARX1 \regf_reg[30][30]  ( .D(n1037), .CLK(clk), .RSTB(n2623), .Q(
        \regf[30][30] ) );
  DFFARX1 \regf_reg[30][29]  ( .D(n1036), .CLK(clk), .RSTB(n2623), .Q(
        \regf[30][29] ) );
  DFFARX1 \regf_reg[30][28]  ( .D(n1035), .CLK(clk), .RSTB(n2623), .Q(
        \regf[30][28] ) );
  DFFARX1 \regf_reg[30][27]  ( .D(n1034), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][27] ) );
  DFFARX1 \regf_reg[30][26]  ( .D(n1033), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][26] ) );
  DFFARX1 \regf_reg[30][25]  ( .D(n1032), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][25] ) );
  DFFARX1 \regf_reg[30][24]  ( .D(n1031), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][24] ) );
  DFFARX1 \regf_reg[30][23]  ( .D(n1030), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][23] ) );
  DFFARX1 \regf_reg[30][22]  ( .D(n1029), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][22] ) );
  DFFARX1 \regf_reg[30][21]  ( .D(n1028), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][21] ) );
  DFFARX1 \regf_reg[30][20]  ( .D(n1027), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][20] ) );
  DFFARX1 \regf_reg[30][19]  ( .D(n1026), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][19] ) );
  DFFARX1 \regf_reg[30][18]  ( .D(n1025), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][18] ) );
  DFFARX1 \regf_reg[30][17]  ( .D(n1024), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][17] ) );
  DFFARX1 \regf_reg[30][16]  ( .D(n1023), .CLK(clk), .RSTB(n2624), .Q(
        \regf[30][16] ) );
  DFFARX1 \regf_reg[30][15]  ( .D(n1022), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][15] ) );
  DFFARX1 \regf_reg[30][14]  ( .D(n1021), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][14] ) );
  DFFARX1 \regf_reg[30][13]  ( .D(n1020), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][13] ) );
  DFFARX1 \regf_reg[30][12]  ( .D(n1019), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][12] ) );
  DFFARX1 \regf_reg[30][11]  ( .D(n1018), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][11] ) );
  DFFARX1 \regf_reg[30][10]  ( .D(n1017), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][10] ) );
  DFFARX1 \regf_reg[30][9]  ( .D(n1016), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][9] ) );
  DFFARX1 \regf_reg[30][8]  ( .D(n1015), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][8] ) );
  DFFARX1 \regf_reg[30][7]  ( .D(n1014), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][7] ) );
  DFFARX1 \regf_reg[30][6]  ( .D(n1013), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][6] ) );
  DFFARX1 \regf_reg[30][5]  ( .D(n1012), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][5] ) );
  DFFARX1 \regf_reg[30][4]  ( .D(n1011), .CLK(clk), .RSTB(n2625), .Q(
        \regf[30][4] ) );
  DFFARX1 \regf_reg[30][3]  ( .D(n1010), .CLK(clk), .RSTB(n2626), .Q(
        \regf[30][3] ) );
  DFFARX1 \regf_reg[30][2]  ( .D(n1009), .CLK(clk), .RSTB(n2626), .Q(
        \regf[30][2] ) );
  DFFARX1 \regf_reg[30][1]  ( .D(n1008), .CLK(clk), .RSTB(n2626), .Q(
        \regf[30][1] ) );
  DFFARX1 \regf_reg[30][0]  ( .D(n1007), .CLK(clk), .RSTB(n2626), .Q(
        \regf[30][0] ) );
  DFFARX1 \regf_reg[29][31]  ( .D(n1006), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][31] ) );
  DFFARX1 \regf_reg[29][30]  ( .D(n1005), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][30] ) );
  DFFARX1 \regf_reg[29][29]  ( .D(n1004), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][29] ) );
  DFFARX1 \regf_reg[29][28]  ( .D(n1003), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][28] ) );
  DFFARX1 \regf_reg[29][27]  ( .D(n1002), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][27] ) );
  DFFARX1 \regf_reg[29][26]  ( .D(n1001), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][26] ) );
  DFFARX1 \regf_reg[29][25]  ( .D(n1000), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][25] ) );
  DFFARX1 \regf_reg[29][24]  ( .D(n999), .CLK(clk), .RSTB(n2626), .Q(
        \regf[29][24] ) );
  DFFARX1 \regf_reg[29][23]  ( .D(n998), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][23] ) );
  DFFARX1 \regf_reg[29][22]  ( .D(n997), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][22] ) );
  DFFARX1 \regf_reg[29][21]  ( .D(n996), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][21] ) );
  DFFARX1 \regf_reg[29][20]  ( .D(n995), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][20] ) );
  DFFARX1 \regf_reg[29][19]  ( .D(n994), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][19] ) );
  DFFARX1 \regf_reg[29][18]  ( .D(n993), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][18] ) );
  DFFARX1 \regf_reg[29][17]  ( .D(n992), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][17] ) );
  DFFARX1 \regf_reg[29][16]  ( .D(n991), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][16] ) );
  DFFARX1 \regf_reg[29][15]  ( .D(n990), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][15] ) );
  DFFARX1 \regf_reg[29][14]  ( .D(n989), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][14] ) );
  DFFARX1 \regf_reg[29][13]  ( .D(n988), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][13] ) );
  DFFARX1 \regf_reg[29][12]  ( .D(n987), .CLK(clk), .RSTB(n2627), .Q(
        \regf[29][12] ) );
  DFFARX1 \regf_reg[29][11]  ( .D(n986), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][11] ) );
  DFFARX1 \regf_reg[29][10]  ( .D(n985), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][10] ) );
  DFFARX1 \regf_reg[29][9]  ( .D(n984), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][9] ) );
  DFFARX1 \regf_reg[29][8]  ( .D(n983), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][8] ) );
  DFFARX1 \regf_reg[29][7]  ( .D(n982), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][7] ) );
  DFFARX1 \regf_reg[29][6]  ( .D(n981), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][6] ) );
  DFFARX1 \regf_reg[29][5]  ( .D(n980), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][5] ) );
  DFFARX1 \regf_reg[29][4]  ( .D(n979), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][4] ) );
  DFFARX1 \regf_reg[29][3]  ( .D(n978), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][3] ) );
  DFFARX1 \regf_reg[29][2]  ( .D(n977), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][2] ) );
  DFFARX1 \regf_reg[29][1]  ( .D(n976), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][1] ) );
  DFFARX1 \regf_reg[29][0]  ( .D(n975), .CLK(clk), .RSTB(n2628), .Q(
        \regf[29][0] ) );
  DFFARX1 \regf_reg[28][31]  ( .D(n974), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][31] ) );
  DFFARX1 \regf_reg[28][30]  ( .D(n973), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][30] ) );
  DFFARX1 \regf_reg[28][29]  ( .D(n972), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][29] ) );
  DFFARX1 \regf_reg[28][28]  ( .D(n971), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][28] ) );
  DFFARX1 \regf_reg[28][27]  ( .D(n970), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][27] ) );
  DFFARX1 \regf_reg[28][26]  ( .D(n969), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][26] ) );
  DFFARX1 \regf_reg[28][25]  ( .D(n968), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][25] ) );
  DFFARX1 \regf_reg[28][24]  ( .D(n967), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][24] ) );
  DFFARX1 \regf_reg[28][23]  ( .D(n966), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][23] ) );
  DFFARX1 \regf_reg[28][22]  ( .D(n965), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][22] ) );
  DFFARX1 \regf_reg[28][21]  ( .D(n964), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][21] ) );
  DFFARX1 \regf_reg[28][20]  ( .D(n963), .CLK(clk), .RSTB(n2629), .Q(
        \regf[28][20] ) );
  DFFARX1 \regf_reg[28][19]  ( .D(n962), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][19] ) );
  DFFARX1 \regf_reg[28][18]  ( .D(n961), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][18] ) );
  DFFARX1 \regf_reg[28][17]  ( .D(n960), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][17] ) );
  DFFARX1 \regf_reg[28][16]  ( .D(n959), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][16] ) );
  DFFARX1 \regf_reg[28][15]  ( .D(n958), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][15] ) );
  DFFARX1 \regf_reg[28][14]  ( .D(n957), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][14] ) );
  DFFARX1 \regf_reg[28][13]  ( .D(n956), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][13] ) );
  DFFARX1 \regf_reg[28][12]  ( .D(n955), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][12] ) );
  DFFARX1 \regf_reg[28][11]  ( .D(n954), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][11] ) );
  DFFARX1 \regf_reg[28][10]  ( .D(n953), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][10] ) );
  DFFARX1 \regf_reg[28][9]  ( .D(n952), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][9] ) );
  DFFARX1 \regf_reg[28][8]  ( .D(n951), .CLK(clk), .RSTB(n2630), .Q(
        \regf[28][8] ) );
  DFFARX1 \regf_reg[28][7]  ( .D(n950), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][7] ) );
  DFFARX1 \regf_reg[28][6]  ( .D(n949), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][6] ) );
  DFFARX1 \regf_reg[28][5]  ( .D(n948), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][5] ) );
  DFFARX1 \regf_reg[28][4]  ( .D(n947), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][4] ) );
  DFFARX1 \regf_reg[28][3]  ( .D(n946), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][3] ) );
  DFFARX1 \regf_reg[28][2]  ( .D(n945), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][2] ) );
  DFFARX1 \regf_reg[28][1]  ( .D(n944), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][1] ) );
  DFFARX1 \regf_reg[28][0]  ( .D(n943), .CLK(clk), .RSTB(n2631), .Q(
        \regf[28][0] ) );
  DFFARX1 \regf_reg[27][31]  ( .D(n942), .CLK(clk), .RSTB(n2631), .Q(
        \regf[27][31] ) );
  DFFARX1 \regf_reg[27][30]  ( .D(n941), .CLK(clk), .RSTB(n2631), .Q(
        \regf[27][30] ) );
  DFFARX1 \regf_reg[27][29]  ( .D(n940), .CLK(clk), .RSTB(n2631), .Q(
        \regf[27][29] ) );
  DFFARX1 \regf_reg[27][28]  ( .D(n939), .CLK(clk), .RSTB(n2631), .Q(
        \regf[27][28] ) );
  DFFARX1 \regf_reg[27][27]  ( .D(n938), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][27] ) );
  DFFARX1 \regf_reg[27][26]  ( .D(n937), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][26] ) );
  DFFARX1 \regf_reg[27][25]  ( .D(n936), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][25] ) );
  DFFARX1 \regf_reg[27][24]  ( .D(n935), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][24] ) );
  DFFARX1 \regf_reg[27][23]  ( .D(n934), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][23] ) );
  DFFARX1 \regf_reg[27][22]  ( .D(n933), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][22] ) );
  DFFARX1 \regf_reg[27][21]  ( .D(n932), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][21] ) );
  DFFARX1 \regf_reg[27][20]  ( .D(n931), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][20] ) );
  DFFARX1 \regf_reg[27][19]  ( .D(n930), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][19] ) );
  DFFARX1 \regf_reg[27][18]  ( .D(n929), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][18] ) );
  DFFARX1 \regf_reg[27][17]  ( .D(n928), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][17] ) );
  DFFARX1 \regf_reg[27][16]  ( .D(n927), .CLK(clk), .RSTB(n2632), .Q(
        \regf[27][16] ) );
  DFFARX1 \regf_reg[27][15]  ( .D(n926), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][15] ) );
  DFFARX1 \regf_reg[27][14]  ( .D(n925), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][14] ) );
  DFFARX1 \regf_reg[27][13]  ( .D(n924), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][13] ) );
  DFFARX1 \regf_reg[27][12]  ( .D(n923), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][12] ) );
  DFFARX1 \regf_reg[27][11]  ( .D(n922), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][11] ) );
  DFFARX1 \regf_reg[27][10]  ( .D(n921), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][10] ) );
  DFFARX1 \regf_reg[27][9]  ( .D(n920), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][9] ) );
  DFFARX1 \regf_reg[27][8]  ( .D(n919), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][8] ) );
  DFFARX1 \regf_reg[27][7]  ( .D(n918), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][7] ) );
  DFFARX1 \regf_reg[27][6]  ( .D(n917), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][6] ) );
  DFFARX1 \regf_reg[27][5]  ( .D(n916), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][5] ) );
  DFFARX1 \regf_reg[27][4]  ( .D(n915), .CLK(clk), .RSTB(n2633), .Q(
        \regf[27][4] ) );
  DFFARX1 \regf_reg[27][3]  ( .D(n914), .CLK(clk), .RSTB(n2634), .Q(
        \regf[27][3] ) );
  DFFARX1 \regf_reg[27][2]  ( .D(n913), .CLK(clk), .RSTB(n2634), .Q(
        \regf[27][2] ) );
  DFFARX1 \regf_reg[27][1]  ( .D(n912), .CLK(clk), .RSTB(n2634), .Q(
        \regf[27][1] ) );
  DFFARX1 \regf_reg[27][0]  ( .D(n911), .CLK(clk), .RSTB(n2634), .Q(
        \regf[27][0] ) );
  DFFARX1 \regf_reg[26][31]  ( .D(n910), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][31] ) );
  DFFARX1 \regf_reg[26][30]  ( .D(n909), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][30] ) );
  DFFARX1 \regf_reg[26][29]  ( .D(n908), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][29] ) );
  DFFARX1 \regf_reg[26][28]  ( .D(n907), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][28] ) );
  DFFARX1 \regf_reg[26][27]  ( .D(n906), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][27] ) );
  DFFARX1 \regf_reg[26][26]  ( .D(n905), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][26] ) );
  DFFARX1 \regf_reg[26][25]  ( .D(n904), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][25] ) );
  DFFARX1 \regf_reg[26][24]  ( .D(n903), .CLK(clk), .RSTB(n2634), .Q(
        \regf[26][24] ) );
  DFFARX1 \regf_reg[26][23]  ( .D(n902), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][23] ) );
  DFFARX1 \regf_reg[26][22]  ( .D(n901), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][22] ) );
  DFFARX1 \regf_reg[26][21]  ( .D(n900), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][21] ) );
  DFFARX1 \regf_reg[26][20]  ( .D(n899), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][20] ) );
  DFFARX1 \regf_reg[26][19]  ( .D(n898), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][19] ) );
  DFFARX1 \regf_reg[26][18]  ( .D(n897), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][18] ) );
  DFFARX1 \regf_reg[26][17]  ( .D(n896), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][17] ) );
  DFFARX1 \regf_reg[26][16]  ( .D(n895), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][16] ) );
  DFFARX1 \regf_reg[26][15]  ( .D(n894), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][15] ) );
  DFFARX1 \regf_reg[26][14]  ( .D(n893), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][14] ) );
  DFFARX1 \regf_reg[26][13]  ( .D(n892), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][13] ) );
  DFFARX1 \regf_reg[26][12]  ( .D(n891), .CLK(clk), .RSTB(n2635), .Q(
        \regf[26][12] ) );
  DFFARX1 \regf_reg[26][11]  ( .D(n890), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][11] ) );
  DFFARX1 \regf_reg[26][10]  ( .D(n889), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][10] ) );
  DFFARX1 \regf_reg[26][9]  ( .D(n888), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][9] ) );
  DFFARX1 \regf_reg[26][8]  ( .D(n887), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][8] ) );
  DFFARX1 \regf_reg[26][7]  ( .D(n886), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][7] ) );
  DFFARX1 \regf_reg[26][6]  ( .D(n885), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][6] ) );
  DFFARX1 \regf_reg[26][5]  ( .D(n884), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][5] ) );
  DFFARX1 \regf_reg[26][4]  ( .D(n883), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][4] ) );
  DFFARX1 \regf_reg[26][3]  ( .D(n882), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][3] ) );
  DFFARX1 \regf_reg[26][2]  ( .D(n881), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][2] ) );
  DFFARX1 \regf_reg[26][1]  ( .D(n880), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][1] ) );
  DFFARX1 \regf_reg[26][0]  ( .D(n879), .CLK(clk), .RSTB(n2636), .Q(
        \regf[26][0] ) );
  DFFARX1 \regf_reg[25][31]  ( .D(n878), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][31] ) );
  DFFARX1 \regf_reg[25][30]  ( .D(n877), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][30] ) );
  DFFARX1 \regf_reg[25][29]  ( .D(n876), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][29] ) );
  DFFARX1 \regf_reg[25][28]  ( .D(n875), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][28] ) );
  DFFARX1 \regf_reg[25][27]  ( .D(n874), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][27] ) );
  DFFARX1 \regf_reg[25][26]  ( .D(n873), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][26] ) );
  DFFARX1 \regf_reg[25][25]  ( .D(n872), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][25] ) );
  DFFARX1 \regf_reg[25][24]  ( .D(n871), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][24] ) );
  DFFARX1 \regf_reg[25][23]  ( .D(n870), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][23] ) );
  DFFARX1 \regf_reg[25][22]  ( .D(n869), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][22] ) );
  DFFARX1 \regf_reg[25][21]  ( .D(n868), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][21] ) );
  DFFARX1 \regf_reg[25][20]  ( .D(n867), .CLK(clk), .RSTB(n2637), .Q(
        \regf[25][20] ) );
  DFFARX1 \regf_reg[25][19]  ( .D(n866), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][19] ) );
  DFFARX1 \regf_reg[25][18]  ( .D(n865), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][18] ) );
  DFFARX1 \regf_reg[25][17]  ( .D(n864), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][17] ) );
  DFFARX1 \regf_reg[25][16]  ( .D(n863), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][16] ) );
  DFFARX1 \regf_reg[25][15]  ( .D(n862), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][15] ) );
  DFFARX1 \regf_reg[25][14]  ( .D(n861), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][14] ) );
  DFFARX1 \regf_reg[25][13]  ( .D(n860), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][13] ) );
  DFFARX1 \regf_reg[25][12]  ( .D(n859), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][12] ) );
  DFFARX1 \regf_reg[25][11]  ( .D(n858), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][11] ) );
  DFFARX1 \regf_reg[25][10]  ( .D(n857), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][10] ) );
  DFFARX1 \regf_reg[25][9]  ( .D(n856), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][9] ) );
  DFFARX1 \regf_reg[25][8]  ( .D(n855), .CLK(clk), .RSTB(n2638), .Q(
        \regf[25][8] ) );
  DFFARX1 \regf_reg[25][7]  ( .D(n854), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][7] ) );
  DFFARX1 \regf_reg[25][6]  ( .D(n853), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][6] ) );
  DFFARX1 \regf_reg[25][5]  ( .D(n852), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][5] ) );
  DFFARX1 \regf_reg[25][4]  ( .D(n851), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][4] ) );
  DFFARX1 \regf_reg[25][3]  ( .D(n850), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][3] ) );
  DFFARX1 \regf_reg[25][2]  ( .D(n849), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][2] ) );
  DFFARX1 \regf_reg[25][1]  ( .D(n848), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][1] ) );
  DFFARX1 \regf_reg[25][0]  ( .D(n847), .CLK(clk), .RSTB(n2639), .Q(
        \regf[25][0] ) );
  DFFARX1 \regf_reg[24][31]  ( .D(n846), .CLK(clk), .RSTB(n2639), .Q(
        \regf[24][31] ) );
  DFFARX1 \regf_reg[24][30]  ( .D(n845), .CLK(clk), .RSTB(n2639), .Q(
        \regf[24][30] ) );
  DFFARX1 \regf_reg[24][29]  ( .D(n844), .CLK(clk), .RSTB(n2639), .Q(
        \regf[24][29] ) );
  DFFARX1 \regf_reg[24][28]  ( .D(n843), .CLK(clk), .RSTB(n2639), .Q(
        \regf[24][28] ) );
  DFFARX1 \regf_reg[24][27]  ( .D(n842), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][27] ) );
  DFFARX1 \regf_reg[24][26]  ( .D(n841), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][26] ) );
  DFFARX1 \regf_reg[24][25]  ( .D(n840), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][25] ) );
  DFFARX1 \regf_reg[24][24]  ( .D(n839), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][24] ) );
  DFFARX1 \regf_reg[24][23]  ( .D(n838), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][23] ) );
  DFFARX1 \regf_reg[24][22]  ( .D(n837), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][22] ) );
  DFFARX1 \regf_reg[24][21]  ( .D(n836), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][21] ) );
  DFFARX1 \regf_reg[24][20]  ( .D(n835), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][20] ) );
  DFFARX1 \regf_reg[24][19]  ( .D(n834), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][19] ) );
  DFFARX1 \regf_reg[24][18]  ( .D(n833), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][18] ) );
  DFFARX1 \regf_reg[24][17]  ( .D(n832), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][17] ) );
  DFFARX1 \regf_reg[24][16]  ( .D(n831), .CLK(clk), .RSTB(n2640), .Q(
        \regf[24][16] ) );
  DFFARX1 \regf_reg[24][15]  ( .D(n830), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][15] ) );
  DFFARX1 \regf_reg[24][14]  ( .D(n829), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][14] ) );
  DFFARX1 \regf_reg[24][13]  ( .D(n828), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][13] ) );
  DFFARX1 \regf_reg[24][12]  ( .D(n827), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][12] ) );
  DFFARX1 \regf_reg[24][11]  ( .D(n826), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][11] ) );
  DFFARX1 \regf_reg[24][10]  ( .D(n825), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][10] ) );
  DFFARX1 \regf_reg[24][9]  ( .D(n824), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][9] ) );
  DFFARX1 \regf_reg[24][8]  ( .D(n823), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][8] ) );
  DFFARX1 \regf_reg[24][7]  ( .D(n822), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][7] ) );
  DFFARX1 \regf_reg[24][6]  ( .D(n821), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][6] ) );
  DFFARX1 \regf_reg[24][5]  ( .D(n820), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][5] ) );
  DFFARX1 \regf_reg[24][4]  ( .D(n819), .CLK(clk), .RSTB(n2641), .Q(
        \regf[24][4] ) );
  DFFARX1 \regf_reg[24][3]  ( .D(n818), .CLK(clk), .RSTB(n2642), .Q(
        \regf[24][3] ) );
  DFFARX1 \regf_reg[24][2]  ( .D(n817), .CLK(clk), .RSTB(n2642), .Q(
        \regf[24][2] ) );
  DFFARX1 \regf_reg[24][1]  ( .D(n816), .CLK(clk), .RSTB(n2642), .Q(
        \regf[24][1] ) );
  DFFARX1 \regf_reg[24][0]  ( .D(n815), .CLK(clk), .RSTB(n2642), .Q(
        \regf[24][0] ) );
  DFFARX1 \regf_reg[23][31]  ( .D(n814), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][31] ) );
  DFFARX1 \regf_reg[23][30]  ( .D(n813), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][30] ) );
  DFFARX1 \regf_reg[23][29]  ( .D(n812), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][29] ) );
  DFFARX1 \regf_reg[23][28]  ( .D(n811), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][28] ) );
  DFFARX1 \regf_reg[23][27]  ( .D(n810), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][27] ) );
  DFFARX1 \regf_reg[23][26]  ( .D(n809), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][26] ) );
  DFFARX1 \regf_reg[23][25]  ( .D(n808), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][25] ) );
  DFFARX1 \regf_reg[23][24]  ( .D(n807), .CLK(clk), .RSTB(n2642), .Q(
        \regf[23][24] ) );
  DFFARX1 \regf_reg[23][23]  ( .D(n806), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][23] ) );
  DFFARX1 \regf_reg[23][22]  ( .D(n805), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][22] ) );
  DFFARX1 \regf_reg[23][21]  ( .D(n804), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][21] ) );
  DFFARX1 \regf_reg[23][20]  ( .D(n803), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][20] ) );
  DFFARX1 \regf_reg[23][19]  ( .D(n802), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][19] ) );
  DFFARX1 \regf_reg[23][18]  ( .D(n801), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][18] ) );
  DFFARX1 \regf_reg[23][17]  ( .D(n800), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][17] ) );
  DFFARX1 \regf_reg[23][16]  ( .D(n799), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][16] ) );
  DFFARX1 \regf_reg[23][15]  ( .D(n798), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][15] ) );
  DFFARX1 \regf_reg[23][14]  ( .D(n797), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][14] ) );
  DFFARX1 \regf_reg[23][13]  ( .D(n796), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][13] ) );
  DFFARX1 \regf_reg[23][12]  ( .D(n795), .CLK(clk), .RSTB(n2643), .Q(
        \regf[23][12] ) );
  DFFARX1 \regf_reg[23][11]  ( .D(n794), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][11] ) );
  DFFARX1 \regf_reg[23][10]  ( .D(n793), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][10] ) );
  DFFARX1 \regf_reg[23][9]  ( .D(n792), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][9] ) );
  DFFARX1 \regf_reg[23][8]  ( .D(n791), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][8] ) );
  DFFARX1 \regf_reg[23][7]  ( .D(n790), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][7] ) );
  DFFARX1 \regf_reg[23][6]  ( .D(n789), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][6] ) );
  DFFARX1 \regf_reg[23][5]  ( .D(n788), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][5] ) );
  DFFARX1 \regf_reg[23][4]  ( .D(n787), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][4] ) );
  DFFARX1 \regf_reg[23][3]  ( .D(n786), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][3] ) );
  DFFARX1 \regf_reg[23][2]  ( .D(n785), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][2] ) );
  DFFARX1 \regf_reg[23][1]  ( .D(n784), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][1] ) );
  DFFARX1 \regf_reg[23][0]  ( .D(n783), .CLK(clk), .RSTB(n2644), .Q(
        \regf[23][0] ) );
  DFFARX1 \regf_reg[22][31]  ( .D(n782), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][31] ) );
  DFFARX1 \regf_reg[22][30]  ( .D(n781), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][30] ) );
  DFFARX1 \regf_reg[22][29]  ( .D(n780), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][29] ) );
  DFFARX1 \regf_reg[22][28]  ( .D(n779), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][28] ) );
  DFFARX1 \regf_reg[22][27]  ( .D(n778), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][27] ) );
  DFFARX1 \regf_reg[22][26]  ( .D(n777), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][26] ) );
  DFFARX1 \regf_reg[22][25]  ( .D(n776), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][25] ) );
  DFFARX1 \regf_reg[22][24]  ( .D(n775), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][24] ) );
  DFFARX1 \regf_reg[22][23]  ( .D(n774), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][23] ) );
  DFFARX1 \regf_reg[22][22]  ( .D(n773), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][22] ) );
  DFFARX1 \regf_reg[22][21]  ( .D(n772), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][21] ) );
  DFFARX1 \regf_reg[22][20]  ( .D(n771), .CLK(clk), .RSTB(n2645), .Q(
        \regf[22][20] ) );
  DFFARX1 \regf_reg[22][19]  ( .D(n770), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][19] ) );
  DFFARX1 \regf_reg[22][18]  ( .D(n769), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][18] ) );
  DFFARX1 \regf_reg[22][17]  ( .D(n768), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][17] ) );
  DFFARX1 \regf_reg[22][16]  ( .D(n767), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][16] ) );
  DFFARX1 \regf_reg[22][15]  ( .D(n766), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][15] ) );
  DFFARX1 \regf_reg[22][14]  ( .D(n765), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][14] ) );
  DFFARX1 \regf_reg[22][13]  ( .D(n764), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][13] ) );
  DFFARX1 \regf_reg[22][12]  ( .D(n763), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][12] ) );
  DFFARX1 \regf_reg[22][11]  ( .D(n762), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][11] ) );
  DFFARX1 \regf_reg[22][10]  ( .D(n761), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][10] ) );
  DFFARX1 \regf_reg[22][9]  ( .D(n760), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][9] ) );
  DFFARX1 \regf_reg[22][8]  ( .D(n759), .CLK(clk), .RSTB(n2646), .Q(
        \regf[22][8] ) );
  DFFARX1 \regf_reg[22][7]  ( .D(n758), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][7] ) );
  DFFARX1 \regf_reg[22][6]  ( .D(n757), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][6] ) );
  DFFARX1 \regf_reg[22][5]  ( .D(n756), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][5] ) );
  DFFARX1 \regf_reg[22][4]  ( .D(n755), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][4] ) );
  DFFARX1 \regf_reg[22][3]  ( .D(n754), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][3] ) );
  DFFARX1 \regf_reg[22][2]  ( .D(n753), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][2] ) );
  DFFARX1 \regf_reg[22][1]  ( .D(n752), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][1] ) );
  DFFARX1 \regf_reg[22][0]  ( .D(n751), .CLK(clk), .RSTB(n2647), .Q(
        \regf[22][0] ) );
  DFFARX1 \regf_reg[21][31]  ( .D(n750), .CLK(clk), .RSTB(n2647), .Q(
        \regf[21][31] ) );
  DFFARX1 \regf_reg[21][30]  ( .D(n749), .CLK(clk), .RSTB(n2647), .Q(
        \regf[21][30] ) );
  DFFARX1 \regf_reg[21][29]  ( .D(n748), .CLK(clk), .RSTB(n2647), .Q(
        \regf[21][29] ) );
  DFFARX1 \regf_reg[21][28]  ( .D(n747), .CLK(clk), .RSTB(n2647), .Q(
        \regf[21][28] ) );
  DFFARX1 \regf_reg[21][27]  ( .D(n746), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][27] ) );
  DFFARX1 \regf_reg[21][26]  ( .D(n745), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][26] ) );
  DFFARX1 \regf_reg[21][25]  ( .D(n744), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][25] ) );
  DFFARX1 \regf_reg[21][24]  ( .D(n743), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][24] ) );
  DFFARX1 \regf_reg[21][23]  ( .D(n742), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][23] ) );
  DFFARX1 \regf_reg[21][22]  ( .D(n741), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][22] ) );
  DFFARX1 \regf_reg[21][21]  ( .D(n740), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][21] ) );
  DFFARX1 \regf_reg[21][20]  ( .D(n739), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][20] ) );
  DFFARX1 \regf_reg[21][19]  ( .D(n738), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][19] ) );
  DFFARX1 \regf_reg[21][18]  ( .D(n737), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][18] ) );
  DFFARX1 \regf_reg[21][17]  ( .D(n736), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][17] ) );
  DFFARX1 \regf_reg[21][16]  ( .D(n735), .CLK(clk), .RSTB(n2648), .Q(
        \regf[21][16] ) );
  DFFARX1 \regf_reg[21][15]  ( .D(n734), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][15] ) );
  DFFARX1 \regf_reg[21][14]  ( .D(n733), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][14] ) );
  DFFARX1 \regf_reg[21][13]  ( .D(n732), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][13] ) );
  DFFARX1 \regf_reg[21][12]  ( .D(n731), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][12] ) );
  DFFARX1 \regf_reg[21][11]  ( .D(n730), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][11] ) );
  DFFARX1 \regf_reg[21][10]  ( .D(n729), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][10] ) );
  DFFARX1 \regf_reg[21][9]  ( .D(n728), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][9] ) );
  DFFARX1 \regf_reg[21][8]  ( .D(n727), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][8] ) );
  DFFARX1 \regf_reg[21][7]  ( .D(n726), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][7] ) );
  DFFARX1 \regf_reg[21][6]  ( .D(n725), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][6] ) );
  DFFARX1 \regf_reg[21][5]  ( .D(n724), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][5] ) );
  DFFARX1 \regf_reg[21][4]  ( .D(n723), .CLK(clk), .RSTB(n2649), .Q(
        \regf[21][4] ) );
  DFFARX1 \regf_reg[21][3]  ( .D(n722), .CLK(clk), .RSTB(n2650), .Q(
        \regf[21][3] ) );
  DFFARX1 \regf_reg[21][2]  ( .D(n721), .CLK(clk), .RSTB(n2650), .Q(
        \regf[21][2] ) );
  DFFARX1 \regf_reg[21][1]  ( .D(n720), .CLK(clk), .RSTB(n2650), .Q(
        \regf[21][1] ) );
  DFFARX1 \regf_reg[21][0]  ( .D(n719), .CLK(clk), .RSTB(n2650), .Q(
        \regf[21][0] ) );
  DFFARX1 \regf_reg[20][31]  ( .D(n718), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][31] ) );
  DFFARX1 \regf_reg[20][30]  ( .D(n717), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][30] ) );
  DFFARX1 \regf_reg[20][29]  ( .D(n716), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][29] ) );
  DFFARX1 \regf_reg[20][28]  ( .D(n715), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][28] ) );
  DFFARX1 \regf_reg[20][27]  ( .D(n714), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][27] ) );
  DFFARX1 \regf_reg[20][26]  ( .D(n713), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][26] ) );
  DFFARX1 \regf_reg[20][25]  ( .D(n712), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][25] ) );
  DFFARX1 \regf_reg[20][24]  ( .D(n711), .CLK(clk), .RSTB(n2650), .Q(
        \regf[20][24] ) );
  DFFARX1 \regf_reg[20][23]  ( .D(n710), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][23] ) );
  DFFARX1 \regf_reg[20][22]  ( .D(n709), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][22] ) );
  DFFARX1 \regf_reg[20][21]  ( .D(n708), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][21] ) );
  DFFARX1 \regf_reg[20][20]  ( .D(n707), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][20] ) );
  DFFARX1 \regf_reg[20][19]  ( .D(n706), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][19] ) );
  DFFARX1 \regf_reg[20][18]  ( .D(n705), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][18] ) );
  DFFARX1 \regf_reg[20][17]  ( .D(n704), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][17] ) );
  DFFARX1 \regf_reg[20][16]  ( .D(n703), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][16] ) );
  DFFARX1 \regf_reg[20][15]  ( .D(n702), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][15] ) );
  DFFARX1 \regf_reg[20][14]  ( .D(n701), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][14] ) );
  DFFARX1 \regf_reg[20][13]  ( .D(n700), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][13] ) );
  DFFARX1 \regf_reg[20][12]  ( .D(n699), .CLK(clk), .RSTB(n2651), .Q(
        \regf[20][12] ) );
  DFFARX1 \regf_reg[20][11]  ( .D(n698), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][11] ) );
  DFFARX1 \regf_reg[20][10]  ( .D(n697), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][10] ) );
  DFFARX1 \regf_reg[20][9]  ( .D(n696), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][9] ) );
  DFFARX1 \regf_reg[20][8]  ( .D(n695), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][8] ) );
  DFFARX1 \regf_reg[20][7]  ( .D(n694), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][7] ) );
  DFFARX1 \regf_reg[20][6]  ( .D(n693), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][6] ) );
  DFFARX1 \regf_reg[20][5]  ( .D(n692), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][5] ) );
  DFFARX1 \regf_reg[20][4]  ( .D(n691), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][4] ) );
  DFFARX1 \regf_reg[20][3]  ( .D(n690), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][3] ) );
  DFFARX1 \regf_reg[20][2]  ( .D(n689), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][2] ) );
  DFFARX1 \regf_reg[20][1]  ( .D(n688), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][1] ) );
  DFFARX1 \regf_reg[20][0]  ( .D(n687), .CLK(clk), .RSTB(n2652), .Q(
        \regf[20][0] ) );
  DFFARX1 \regf_reg[19][31]  ( .D(n686), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][31] ) );
  DFFARX1 \regf_reg[19][30]  ( .D(n685), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][30] ) );
  DFFARX1 \regf_reg[19][29]  ( .D(n684), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][29] ) );
  DFFARX1 \regf_reg[19][28]  ( .D(n683), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][28] ) );
  DFFARX1 \regf_reg[19][27]  ( .D(n682), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][27] ) );
  DFFARX1 \regf_reg[19][26]  ( .D(n681), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][26] ) );
  DFFARX1 \regf_reg[19][25]  ( .D(n680), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][25] ) );
  DFFARX1 \regf_reg[19][24]  ( .D(n679), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][24] ) );
  DFFARX1 \regf_reg[19][23]  ( .D(n678), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][23] ) );
  DFFARX1 \regf_reg[19][22]  ( .D(n677), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][22] ) );
  DFFARX1 \regf_reg[19][21]  ( .D(n676), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][21] ) );
  DFFARX1 \regf_reg[19][20]  ( .D(n675), .CLK(clk), .RSTB(n2653), .Q(
        \regf[19][20] ) );
  DFFARX1 \regf_reg[19][19]  ( .D(n674), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][19] ) );
  DFFARX1 \regf_reg[19][18]  ( .D(n673), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][18] ) );
  DFFARX1 \regf_reg[19][17]  ( .D(n672), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][17] ) );
  DFFARX1 \regf_reg[19][16]  ( .D(n671), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][16] ) );
  DFFARX1 \regf_reg[19][15]  ( .D(n670), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][15] ) );
  DFFARX1 \regf_reg[19][14]  ( .D(n669), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][14] ) );
  DFFARX1 \regf_reg[19][13]  ( .D(n668), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][13] ) );
  DFFARX1 \regf_reg[19][12]  ( .D(n667), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][12] ) );
  DFFARX1 \regf_reg[19][11]  ( .D(n666), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][11] ) );
  DFFARX1 \regf_reg[19][10]  ( .D(n665), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][10] ) );
  DFFARX1 \regf_reg[19][9]  ( .D(n664), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][9] ) );
  DFFARX1 \regf_reg[19][8]  ( .D(n663), .CLK(clk), .RSTB(n2654), .Q(
        \regf[19][8] ) );
  DFFARX1 \regf_reg[19][7]  ( .D(n662), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][7] ) );
  DFFARX1 \regf_reg[19][6]  ( .D(n661), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][6] ) );
  DFFARX1 \regf_reg[19][5]  ( .D(n660), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][5] ) );
  DFFARX1 \regf_reg[19][4]  ( .D(n659), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][4] ) );
  DFFARX1 \regf_reg[19][3]  ( .D(n658), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][3] ) );
  DFFARX1 \regf_reg[19][2]  ( .D(n657), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][2] ) );
  DFFARX1 \regf_reg[19][1]  ( .D(n656), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][1] ) );
  DFFARX1 \regf_reg[19][0]  ( .D(n655), .CLK(clk), .RSTB(n2655), .Q(
        \regf[19][0] ) );
  DFFARX1 \regf_reg[18][31]  ( .D(n654), .CLK(clk), .RSTB(n2655), .Q(
        \regf[18][31] ) );
  DFFARX1 \regf_reg[18][30]  ( .D(n653), .CLK(clk), .RSTB(n2655), .Q(
        \regf[18][30] ) );
  DFFARX1 \regf_reg[18][29]  ( .D(n652), .CLK(clk), .RSTB(n2655), .Q(
        \regf[18][29] ) );
  DFFARX1 \regf_reg[18][28]  ( .D(n651), .CLK(clk), .RSTB(n2655), .Q(
        \regf[18][28] ) );
  DFFARX1 \regf_reg[18][27]  ( .D(n650), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][27] ) );
  DFFARX1 \regf_reg[18][26]  ( .D(n649), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][26] ) );
  DFFARX1 \regf_reg[18][25]  ( .D(n648), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][25] ) );
  DFFARX1 \regf_reg[18][24]  ( .D(n647), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][24] ) );
  DFFARX1 \regf_reg[18][23]  ( .D(n646), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][23] ) );
  DFFARX1 \regf_reg[18][22]  ( .D(n645), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][22] ) );
  DFFARX1 \regf_reg[18][21]  ( .D(n644), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][21] ) );
  DFFARX1 \regf_reg[18][20]  ( .D(n643), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][20] ) );
  DFFARX1 \regf_reg[18][19]  ( .D(n642), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][19] ) );
  DFFARX1 \regf_reg[18][18]  ( .D(n641), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][18] ) );
  DFFARX1 \regf_reg[18][17]  ( .D(n640), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][17] ) );
  DFFARX1 \regf_reg[18][16]  ( .D(n639), .CLK(clk), .RSTB(n2656), .Q(
        \regf[18][16] ) );
  DFFARX1 \regf_reg[18][15]  ( .D(n638), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][15] ) );
  DFFARX1 \regf_reg[18][14]  ( .D(n637), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][14] ) );
  DFFARX1 \regf_reg[18][13]  ( .D(n636), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][13] ) );
  DFFARX1 \regf_reg[18][12]  ( .D(n635), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][12] ) );
  DFFARX1 \regf_reg[18][11]  ( .D(n634), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][11] ) );
  DFFARX1 \regf_reg[18][10]  ( .D(n633), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][10] ) );
  DFFARX1 \regf_reg[18][9]  ( .D(n632), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][9] ) );
  DFFARX1 \regf_reg[18][8]  ( .D(n631), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][8] ) );
  DFFARX1 \regf_reg[18][7]  ( .D(n630), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][7] ) );
  DFFARX1 \regf_reg[18][6]  ( .D(n629), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][6] ) );
  DFFARX1 \regf_reg[18][5]  ( .D(n628), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][5] ) );
  DFFARX1 \regf_reg[18][4]  ( .D(n627), .CLK(clk), .RSTB(n2657), .Q(
        \regf[18][4] ) );
  DFFARX1 \regf_reg[18][3]  ( .D(n626), .CLK(clk), .RSTB(n2658), .Q(
        \regf[18][3] ) );
  DFFARX1 \regf_reg[18][2]  ( .D(n625), .CLK(clk), .RSTB(n2658), .Q(
        \regf[18][2] ) );
  DFFARX1 \regf_reg[18][1]  ( .D(n624), .CLK(clk), .RSTB(n2658), .Q(
        \regf[18][1] ) );
  DFFARX1 \regf_reg[18][0]  ( .D(n623), .CLK(clk), .RSTB(n2658), .Q(
        \regf[18][0] ) );
  DFFARX1 \regf_reg[17][31]  ( .D(n622), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][31] ) );
  DFFARX1 \regf_reg[17][30]  ( .D(n621), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][30] ) );
  DFFARX1 \regf_reg[17][29]  ( .D(n620), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][29] ) );
  DFFARX1 \regf_reg[17][28]  ( .D(n619), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][28] ) );
  DFFARX1 \regf_reg[17][27]  ( .D(n618), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][27] ) );
  DFFARX1 \regf_reg[17][26]  ( .D(n617), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][26] ) );
  DFFARX1 \regf_reg[17][25]  ( .D(n616), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][25] ) );
  DFFARX1 \regf_reg[17][24]  ( .D(n615), .CLK(clk), .RSTB(n2658), .Q(
        \regf[17][24] ) );
  DFFARX1 \regf_reg[17][23]  ( .D(n614), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][23] ) );
  DFFARX1 \regf_reg[17][22]  ( .D(n613), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][22] ) );
  DFFARX1 \regf_reg[17][21]  ( .D(n612), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][21] ) );
  DFFARX1 \regf_reg[17][20]  ( .D(n611), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][20] ) );
  DFFARX1 \regf_reg[17][19]  ( .D(n610), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][19] ) );
  DFFARX1 \regf_reg[17][18]  ( .D(n609), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][18] ) );
  DFFARX1 \regf_reg[17][17]  ( .D(n608), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][17] ) );
  DFFARX1 \regf_reg[17][16]  ( .D(n607), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][16] ) );
  DFFARX1 \regf_reg[17][15]  ( .D(n606), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][15] ) );
  DFFARX1 \regf_reg[17][14]  ( .D(n605), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][14] ) );
  DFFARX1 \regf_reg[17][13]  ( .D(n604), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][13] ) );
  DFFARX1 \regf_reg[17][12]  ( .D(n603), .CLK(clk), .RSTB(n2659), .Q(
        \regf[17][12] ) );
  DFFARX1 \regf_reg[17][11]  ( .D(n602), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][11] ) );
  DFFARX1 \regf_reg[17][10]  ( .D(n601), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][10] ) );
  DFFARX1 \regf_reg[17][9]  ( .D(n600), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][9] ) );
  DFFARX1 \regf_reg[17][8]  ( .D(n599), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][8] ) );
  DFFARX1 \regf_reg[17][7]  ( .D(n598), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][7] ) );
  DFFARX1 \regf_reg[17][6]  ( .D(n597), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][6] ) );
  DFFARX1 \regf_reg[17][5]  ( .D(n596), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][5] ) );
  DFFARX1 \regf_reg[17][4]  ( .D(n595), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][4] ) );
  DFFARX1 \regf_reg[17][3]  ( .D(n594), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][3] ) );
  DFFARX1 \regf_reg[17][2]  ( .D(n593), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][2] ) );
  DFFARX1 \regf_reg[17][1]  ( .D(n592), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][1] ) );
  DFFARX1 \regf_reg[17][0]  ( .D(n591), .CLK(clk), .RSTB(n2660), .Q(
        \regf[17][0] ) );
  DFFARX1 \regf_reg[16][31]  ( .D(n590), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][31] ) );
  DFFARX1 \regf_reg[16][30]  ( .D(n589), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][30] ) );
  DFFARX1 \regf_reg[16][29]  ( .D(n588), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][29] ) );
  DFFARX1 \regf_reg[16][28]  ( .D(n587), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][28] ) );
  DFFARX1 \regf_reg[16][27]  ( .D(n586), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][27] ) );
  DFFARX1 \regf_reg[16][26]  ( .D(n585), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][26] ) );
  DFFARX1 \regf_reg[16][25]  ( .D(n584), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][25] ) );
  DFFARX1 \regf_reg[16][24]  ( .D(n583), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][24] ) );
  DFFARX1 \regf_reg[16][23]  ( .D(n582), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][23] ) );
  DFFARX1 \regf_reg[16][22]  ( .D(n581), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][22] ) );
  DFFARX1 \regf_reg[16][21]  ( .D(n580), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][21] ) );
  DFFARX1 \regf_reg[16][20]  ( .D(n579), .CLK(clk), .RSTB(n2661), .Q(
        \regf[16][20] ) );
  DFFARX1 \regf_reg[16][19]  ( .D(n578), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][19] ) );
  DFFARX1 \regf_reg[16][18]  ( .D(n577), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][18] ) );
  DFFARX1 \regf_reg[16][17]  ( .D(n576), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][17] ) );
  DFFARX1 \regf_reg[16][16]  ( .D(n575), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][16] ) );
  DFFARX1 \regf_reg[16][15]  ( .D(n574), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][15] ) );
  DFFARX1 \regf_reg[16][14]  ( .D(n573), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][14] ) );
  DFFARX1 \regf_reg[16][13]  ( .D(n572), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][13] ) );
  DFFARX1 \regf_reg[16][12]  ( .D(n571), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][12] ) );
  DFFARX1 \regf_reg[16][11]  ( .D(n570), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][11] ) );
  DFFARX1 \regf_reg[16][10]  ( .D(n569), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][10] ) );
  DFFARX1 \regf_reg[16][9]  ( .D(n568), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][9] ) );
  DFFARX1 \regf_reg[16][8]  ( .D(n567), .CLK(clk), .RSTB(n2662), .Q(
        \regf[16][8] ) );
  DFFARX1 \regf_reg[16][7]  ( .D(n566), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][7] ) );
  DFFARX1 \regf_reg[16][6]  ( .D(n565), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][6] ) );
  DFFARX1 \regf_reg[16][5]  ( .D(n564), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][5] ) );
  DFFARX1 \regf_reg[16][4]  ( .D(n563), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][4] ) );
  DFFARX1 \regf_reg[16][3]  ( .D(n562), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][3] ) );
  DFFARX1 \regf_reg[16][2]  ( .D(n561), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][2] ) );
  DFFARX1 \regf_reg[16][1]  ( .D(n560), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][1] ) );
  DFFARX1 \regf_reg[16][0]  ( .D(n559), .CLK(clk), .RSTB(n2663), .Q(
        \regf[16][0] ) );
  DFFARX1 \regf_reg[15][31]  ( .D(n558), .CLK(clk), .RSTB(n2663), .Q(
        \regf[15][31] ) );
  DFFARX1 \regf_reg[15][30]  ( .D(n557), .CLK(clk), .RSTB(n2663), .Q(
        \regf[15][30] ) );
  DFFARX1 \regf_reg[15][29]  ( .D(n556), .CLK(clk), .RSTB(n2663), .Q(
        \regf[15][29] ) );
  DFFARX1 \regf_reg[15][28]  ( .D(n555), .CLK(clk), .RSTB(n2663), .Q(
        \regf[15][28] ) );
  DFFARX1 \regf_reg[15][27]  ( .D(n554), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][27] ) );
  DFFARX1 \regf_reg[15][26]  ( .D(n553), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][26] ) );
  DFFARX1 \regf_reg[15][25]  ( .D(n552), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][25] ) );
  DFFARX1 \regf_reg[15][24]  ( .D(n551), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][24] ) );
  DFFARX1 \regf_reg[15][23]  ( .D(n550), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][23] ) );
  DFFARX1 \regf_reg[15][22]  ( .D(n549), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][22] ) );
  DFFARX1 \regf_reg[15][21]  ( .D(n548), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][21] ) );
  DFFARX1 \regf_reg[15][20]  ( .D(n547), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][20] ) );
  DFFARX1 \regf_reg[15][19]  ( .D(n546), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][19] ) );
  DFFARX1 \regf_reg[15][18]  ( .D(n545), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][18] ) );
  DFFARX1 \regf_reg[15][17]  ( .D(n544), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][17] ) );
  DFFARX1 \regf_reg[15][16]  ( .D(n543), .CLK(clk), .RSTB(n2664), .Q(
        \regf[15][16] ) );
  DFFARX1 \regf_reg[15][15]  ( .D(n542), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][15] ) );
  DFFARX1 \regf_reg[15][14]  ( .D(n541), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][14] ) );
  DFFARX1 \regf_reg[15][13]  ( .D(n540), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][13] ) );
  DFFARX1 \regf_reg[15][12]  ( .D(n539), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][12] ) );
  DFFARX1 \regf_reg[15][11]  ( .D(n538), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][11] ) );
  DFFARX1 \regf_reg[15][10]  ( .D(n537), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][10] ) );
  DFFARX1 \regf_reg[15][9]  ( .D(n536), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][9] ) );
  DFFARX1 \regf_reg[15][8]  ( .D(n535), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][8] ) );
  DFFARX1 \regf_reg[15][7]  ( .D(n534), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][7] ) );
  DFFARX1 \regf_reg[15][6]  ( .D(n533), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][6] ) );
  DFFARX1 \regf_reg[15][5]  ( .D(n532), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][5] ) );
  DFFARX1 \regf_reg[15][4]  ( .D(n531), .CLK(clk), .RSTB(n2665), .Q(
        \regf[15][4] ) );
  DFFARX1 \regf_reg[15][3]  ( .D(n530), .CLK(clk), .RSTB(n2666), .Q(
        \regf[15][3] ) );
  DFFARX1 \regf_reg[15][2]  ( .D(n529), .CLK(clk), .RSTB(n2666), .Q(
        \regf[15][2] ) );
  DFFARX1 \regf_reg[15][1]  ( .D(n528), .CLK(clk), .RSTB(n2666), .Q(
        \regf[15][1] ) );
  DFFARX1 \regf_reg[15][0]  ( .D(n527), .CLK(clk), .RSTB(n2666), .Q(
        \regf[15][0] ) );
  DFFARX1 \regf_reg[14][31]  ( .D(n526), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][31] ) );
  DFFARX1 \regf_reg[14][30]  ( .D(n525), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][30] ) );
  DFFARX1 \regf_reg[14][29]  ( .D(n524), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][29] ) );
  DFFARX1 \regf_reg[14][28]  ( .D(n523), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][28] ) );
  DFFARX1 \regf_reg[14][27]  ( .D(n522), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][27] ) );
  DFFARX1 \regf_reg[14][26]  ( .D(n521), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][26] ) );
  DFFARX1 \regf_reg[14][25]  ( .D(n520), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][25] ) );
  DFFARX1 \regf_reg[14][24]  ( .D(n519), .CLK(clk), .RSTB(n2666), .Q(
        \regf[14][24] ) );
  DFFARX1 \regf_reg[14][23]  ( .D(n518), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][23] ) );
  DFFARX1 \regf_reg[14][22]  ( .D(n517), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][22] ) );
  DFFARX1 \regf_reg[14][21]  ( .D(n516), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][21] ) );
  DFFARX1 \regf_reg[14][20]  ( .D(n515), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][20] ) );
  DFFARX1 \regf_reg[14][19]  ( .D(n514), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][19] ) );
  DFFARX1 \regf_reg[14][18]  ( .D(n513), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][18] ) );
  DFFARX1 \regf_reg[14][17]  ( .D(n512), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][17] ) );
  DFFARX1 \regf_reg[14][16]  ( .D(n511), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][16] ) );
  DFFARX1 \regf_reg[14][15]  ( .D(n510), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][15] ) );
  DFFARX1 \regf_reg[14][14]  ( .D(n509), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][14] ) );
  DFFARX1 \regf_reg[14][13]  ( .D(n508), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][13] ) );
  DFFARX1 \regf_reg[14][12]  ( .D(n507), .CLK(clk), .RSTB(n2667), .Q(
        \regf[14][12] ) );
  DFFARX1 \regf_reg[14][11]  ( .D(n506), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][11] ) );
  DFFARX1 \regf_reg[14][10]  ( .D(n505), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][10] ) );
  DFFARX1 \regf_reg[14][9]  ( .D(n504), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][9] ) );
  DFFARX1 \regf_reg[14][8]  ( .D(n503), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][8] ) );
  DFFARX1 \regf_reg[14][7]  ( .D(n502), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][7] ) );
  DFFARX1 \regf_reg[14][6]  ( .D(n501), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][6] ) );
  DFFARX1 \regf_reg[14][5]  ( .D(n500), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][5] ) );
  DFFARX1 \regf_reg[14][4]  ( .D(n499), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][4] ) );
  DFFARX1 \regf_reg[14][3]  ( .D(n498), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][3] ) );
  DFFARX1 \regf_reg[14][2]  ( .D(n497), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][2] ) );
  DFFARX1 \regf_reg[14][1]  ( .D(n496), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][1] ) );
  DFFARX1 \regf_reg[14][0]  ( .D(n495), .CLK(clk), .RSTB(n2668), .Q(
        \regf[14][0] ) );
  DFFARX1 \regf_reg[13][31]  ( .D(n494), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][31] ) );
  DFFARX1 \regf_reg[13][30]  ( .D(n493), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][30] ) );
  DFFARX1 \regf_reg[13][29]  ( .D(n492), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][29] ) );
  DFFARX1 \regf_reg[13][28]  ( .D(n491), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][28] ) );
  DFFARX1 \regf_reg[13][27]  ( .D(n490), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][27] ) );
  DFFARX1 \regf_reg[13][26]  ( .D(n489), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][26] ) );
  DFFARX1 \regf_reg[13][25]  ( .D(n488), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][25] ) );
  DFFARX1 \regf_reg[13][24]  ( .D(n487), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][24] ) );
  DFFARX1 \regf_reg[13][23]  ( .D(n486), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][23] ) );
  DFFARX1 \regf_reg[13][22]  ( .D(n485), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][22] ) );
  DFFARX1 \regf_reg[13][21]  ( .D(n484), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][21] ) );
  DFFARX1 \regf_reg[13][20]  ( .D(n483), .CLK(clk), .RSTB(n2669), .Q(
        \regf[13][20] ) );
  DFFARX1 \regf_reg[13][19]  ( .D(n482), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][19] ) );
  DFFARX1 \regf_reg[13][18]  ( .D(n481), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][18] ) );
  DFFARX1 \regf_reg[13][17]  ( .D(n480), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][17] ) );
  DFFARX1 \regf_reg[13][16]  ( .D(n479), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][16] ) );
  DFFARX1 \regf_reg[13][15]  ( .D(n478), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][15] ) );
  DFFARX1 \regf_reg[13][14]  ( .D(n477), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][14] ) );
  DFFARX1 \regf_reg[13][13]  ( .D(n476), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][13] ) );
  DFFARX1 \regf_reg[13][12]  ( .D(n475), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][12] ) );
  DFFARX1 \regf_reg[13][11]  ( .D(n474), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][11] ) );
  DFFARX1 \regf_reg[13][10]  ( .D(n473), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][10] ) );
  DFFARX1 \regf_reg[13][9]  ( .D(n472), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][9] ) );
  DFFARX1 \regf_reg[13][8]  ( .D(n471), .CLK(clk), .RSTB(n2670), .Q(
        \regf[13][8] ) );
  DFFARX1 \regf_reg[13][7]  ( .D(n470), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][7] ) );
  DFFARX1 \regf_reg[13][6]  ( .D(n469), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][6] ) );
  DFFARX1 \regf_reg[13][5]  ( .D(n468), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][5] ) );
  DFFARX1 \regf_reg[13][4]  ( .D(n467), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][4] ) );
  DFFARX1 \regf_reg[13][3]  ( .D(n466), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][3] ) );
  DFFARX1 \regf_reg[13][2]  ( .D(n465), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][2] ) );
  DFFARX1 \regf_reg[13][1]  ( .D(n464), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][1] ) );
  DFFARX1 \regf_reg[13][0]  ( .D(n463), .CLK(clk), .RSTB(n2671), .Q(
        \regf[13][0] ) );
  DFFARX1 \regf_reg[12][31]  ( .D(n462), .CLK(clk), .RSTB(n2671), .Q(
        \regf[12][31] ) );
  DFFARX1 \regf_reg[12][30]  ( .D(n461), .CLK(clk), .RSTB(n2671), .Q(
        \regf[12][30] ) );
  DFFARX1 \regf_reg[12][29]  ( .D(n460), .CLK(clk), .RSTB(n2671), .Q(
        \regf[12][29] ) );
  DFFARX1 \regf_reg[12][28]  ( .D(n459), .CLK(clk), .RSTB(n2671), .Q(
        \regf[12][28] ) );
  DFFARX1 \regf_reg[12][27]  ( .D(n458), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][27] ) );
  DFFARX1 \regf_reg[12][26]  ( .D(n457), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][26] ) );
  DFFARX1 \regf_reg[12][25]  ( .D(n456), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][25] ) );
  DFFARX1 \regf_reg[12][24]  ( .D(n455), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][24] ) );
  DFFARX1 \regf_reg[12][23]  ( .D(n454), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][23] ) );
  DFFARX1 \regf_reg[12][22]  ( .D(n453), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][22] ) );
  DFFARX1 \regf_reg[12][21]  ( .D(n452), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][21] ) );
  DFFARX1 \regf_reg[12][20]  ( .D(n451), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][20] ) );
  DFFARX1 \regf_reg[12][19]  ( .D(n450), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][19] ) );
  DFFARX1 \regf_reg[12][18]  ( .D(n449), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][18] ) );
  DFFARX1 \regf_reg[12][17]  ( .D(n448), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][17] ) );
  DFFARX1 \regf_reg[12][16]  ( .D(n447), .CLK(clk), .RSTB(n2672), .Q(
        \regf[12][16] ) );
  DFFARX1 \regf_reg[12][15]  ( .D(n446), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][15] ) );
  DFFARX1 \regf_reg[12][14]  ( .D(n445), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][14] ) );
  DFFARX1 \regf_reg[12][13]  ( .D(n444), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][13] ) );
  DFFARX1 \regf_reg[12][12]  ( .D(n443), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][12] ) );
  DFFARX1 \regf_reg[12][11]  ( .D(n442), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][11] ) );
  DFFARX1 \regf_reg[12][10]  ( .D(n441), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][10] ) );
  DFFARX1 \regf_reg[12][9]  ( .D(n440), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][9] ) );
  DFFARX1 \regf_reg[12][8]  ( .D(n439), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][8] ) );
  DFFARX1 \regf_reg[12][7]  ( .D(n438), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][7] ) );
  DFFARX1 \regf_reg[12][6]  ( .D(n437), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][6] ) );
  DFFARX1 \regf_reg[12][5]  ( .D(n436), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][5] ) );
  DFFARX1 \regf_reg[12][4]  ( .D(n435), .CLK(clk), .RSTB(n2673), .Q(
        \regf[12][4] ) );
  DFFARX1 \regf_reg[12][3]  ( .D(n434), .CLK(clk), .RSTB(n2674), .Q(
        \regf[12][3] ) );
  DFFARX1 \regf_reg[12][2]  ( .D(n433), .CLK(clk), .RSTB(n2674), .Q(
        \regf[12][2] ) );
  DFFARX1 \regf_reg[12][1]  ( .D(n432), .CLK(clk), .RSTB(n2674), .Q(
        \regf[12][1] ) );
  DFFARX1 \regf_reg[12][0]  ( .D(n431), .CLK(clk), .RSTB(n2674), .Q(
        \regf[12][0] ) );
  DFFARX1 \regf_reg[11][31]  ( .D(n430), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][31] ) );
  DFFARX1 \regf_reg[11][30]  ( .D(n429), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][30] ) );
  DFFARX1 \regf_reg[11][29]  ( .D(n428), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][29] ) );
  DFFARX1 \regf_reg[11][28]  ( .D(n427), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][28] ) );
  DFFARX1 \regf_reg[11][27]  ( .D(n426), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][27] ) );
  DFFARX1 \regf_reg[11][26]  ( .D(n425), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][26] ) );
  DFFARX1 \regf_reg[11][25]  ( .D(n424), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][25] ) );
  DFFARX1 \regf_reg[11][24]  ( .D(n423), .CLK(clk), .RSTB(n2674), .Q(
        \regf[11][24] ) );
  DFFARX1 \regf_reg[11][23]  ( .D(n422), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][23] ) );
  DFFARX1 \regf_reg[11][22]  ( .D(n421), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][22] ) );
  DFFARX1 \regf_reg[11][21]  ( .D(n420), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][21] ) );
  DFFARX1 \regf_reg[11][20]  ( .D(n419), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][20] ) );
  DFFARX1 \regf_reg[11][19]  ( .D(n418), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][19] ) );
  DFFARX1 \regf_reg[11][18]  ( .D(n417), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][18] ) );
  DFFARX1 \regf_reg[11][17]  ( .D(n416), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][17] ) );
  DFFARX1 \regf_reg[11][16]  ( .D(n415), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][16] ) );
  DFFARX1 \regf_reg[11][15]  ( .D(n414), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][15] ) );
  DFFARX1 \regf_reg[11][14]  ( .D(n413), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][14] ) );
  DFFARX1 \regf_reg[11][13]  ( .D(n412), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][13] ) );
  DFFARX1 \regf_reg[11][12]  ( .D(n411), .CLK(clk), .RSTB(n2675), .Q(
        \regf[11][12] ) );
  DFFARX1 \regf_reg[11][11]  ( .D(n410), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][11] ) );
  DFFARX1 \regf_reg[11][10]  ( .D(n409), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][10] ) );
  DFFARX1 \regf_reg[11][9]  ( .D(n408), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][9] ) );
  DFFARX1 \regf_reg[11][8]  ( .D(n407), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][8] ) );
  DFFARX1 \regf_reg[11][7]  ( .D(n406), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][7] ) );
  DFFARX1 \regf_reg[11][6]  ( .D(n405), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][6] ) );
  DFFARX1 \regf_reg[11][5]  ( .D(n404), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][5] ) );
  DFFARX1 \regf_reg[11][4]  ( .D(n403), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][4] ) );
  DFFARX1 \regf_reg[11][3]  ( .D(n402), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][3] ) );
  DFFARX1 \regf_reg[11][2]  ( .D(n401), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][2] ) );
  DFFARX1 \regf_reg[11][1]  ( .D(n400), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][1] ) );
  DFFARX1 \regf_reg[11][0]  ( .D(n399), .CLK(clk), .RSTB(n2676), .Q(
        \regf[11][0] ) );
  DFFARX1 \regf_reg[10][31]  ( .D(n398), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][31] ) );
  DFFARX1 \regf_reg[10][30]  ( .D(n397), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][30] ) );
  DFFARX1 \regf_reg[10][29]  ( .D(n396), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][29] ) );
  DFFARX1 \regf_reg[10][28]  ( .D(n395), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][28] ) );
  DFFARX1 \regf_reg[10][27]  ( .D(n394), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][27] ) );
  DFFARX1 \regf_reg[10][26]  ( .D(n393), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][26] ) );
  DFFARX1 \regf_reg[10][25]  ( .D(n392), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][25] ) );
  DFFARX1 \regf_reg[10][24]  ( .D(n391), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][24] ) );
  DFFARX1 \regf_reg[10][23]  ( .D(n390), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][23] ) );
  DFFARX1 \regf_reg[10][22]  ( .D(n389), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][22] ) );
  DFFARX1 \regf_reg[10][21]  ( .D(n388), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][21] ) );
  DFFARX1 \regf_reg[10][20]  ( .D(n387), .CLK(clk), .RSTB(n2677), .Q(
        \regf[10][20] ) );
  DFFARX1 \regf_reg[10][19]  ( .D(n386), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][19] ) );
  DFFARX1 \regf_reg[10][18]  ( .D(n385), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][18] ) );
  DFFARX1 \regf_reg[10][17]  ( .D(n384), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][17] ) );
  DFFARX1 \regf_reg[10][16]  ( .D(n383), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][16] ) );
  DFFARX1 \regf_reg[10][15]  ( .D(n382), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][15] ) );
  DFFARX1 \regf_reg[10][14]  ( .D(n381), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][14] ) );
  DFFARX1 \regf_reg[10][13]  ( .D(n380), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][13] ) );
  DFFARX1 \regf_reg[10][12]  ( .D(n379), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][12] ) );
  DFFARX1 \regf_reg[10][11]  ( .D(n378), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][11] ) );
  DFFARX1 \regf_reg[10][10]  ( .D(n377), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][10] ) );
  DFFARX1 \regf_reg[10][9]  ( .D(n376), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][9] ) );
  DFFARX1 \regf_reg[10][8]  ( .D(n375), .CLK(clk), .RSTB(n2678), .Q(
        \regf[10][8] ) );
  DFFARX1 \regf_reg[10][7]  ( .D(n374), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][7] ) );
  DFFARX1 \regf_reg[10][6]  ( .D(n373), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][6] ) );
  DFFARX1 \regf_reg[10][5]  ( .D(n372), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][5] ) );
  DFFARX1 \regf_reg[10][4]  ( .D(n371), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][4] ) );
  DFFARX1 \regf_reg[10][3]  ( .D(n370), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][3] ) );
  DFFARX1 \regf_reg[10][2]  ( .D(n369), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][2] ) );
  DFFARX1 \regf_reg[10][1]  ( .D(n368), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][1] ) );
  DFFARX1 \regf_reg[10][0]  ( .D(n367), .CLK(clk), .RSTB(n2679), .Q(
        \regf[10][0] ) );
  DFFARX1 \regf_reg[9][31]  ( .D(n366), .CLK(clk), .RSTB(n2679), .Q(
        \regf[9][31] ) );
  DFFARX1 \regf_reg[9][30]  ( .D(n365), .CLK(clk), .RSTB(n2679), .Q(
        \regf[9][30] ) );
  DFFARX1 \regf_reg[9][29]  ( .D(n364), .CLK(clk), .RSTB(n2679), .Q(
        \regf[9][29] ) );
  DFFARX1 \regf_reg[9][28]  ( .D(n363), .CLK(clk), .RSTB(n2679), .Q(
        \regf[9][28] ) );
  DFFARX1 \regf_reg[9][27]  ( .D(n362), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][27] ) );
  DFFARX1 \regf_reg[9][26]  ( .D(n361), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][26] ) );
  DFFARX1 \regf_reg[9][25]  ( .D(n360), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][25] ) );
  DFFARX1 \regf_reg[9][24]  ( .D(n359), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][24] ) );
  DFFARX1 \regf_reg[9][23]  ( .D(n358), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][23] ) );
  DFFARX1 \regf_reg[9][22]  ( .D(n357), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][22] ) );
  DFFARX1 \regf_reg[9][21]  ( .D(n356), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][21] ) );
  DFFARX1 \regf_reg[9][20]  ( .D(n355), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][20] ) );
  DFFARX1 \regf_reg[9][19]  ( .D(n354), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][19] ) );
  DFFARX1 \regf_reg[9][18]  ( .D(n353), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][18] ) );
  DFFARX1 \regf_reg[9][17]  ( .D(n352), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][17] ) );
  DFFARX1 \regf_reg[9][16]  ( .D(n351), .CLK(clk), .RSTB(n2680), .Q(
        \regf[9][16] ) );
  DFFARX1 \regf_reg[9][15]  ( .D(n350), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][15] ) );
  DFFARX1 \regf_reg[9][14]  ( .D(n349), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][14] ) );
  DFFARX1 \regf_reg[9][13]  ( .D(n348), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][13] ) );
  DFFARX1 \regf_reg[9][12]  ( .D(n347), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][12] ) );
  DFFARX1 \regf_reg[9][11]  ( .D(n346), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][11] ) );
  DFFARX1 \regf_reg[9][10]  ( .D(n345), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][10] ) );
  DFFARX1 \regf_reg[9][9]  ( .D(n344), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][9] ) );
  DFFARX1 \regf_reg[9][8]  ( .D(n343), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][8] ) );
  DFFARX1 \regf_reg[9][7]  ( .D(n342), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][7] ) );
  DFFARX1 \regf_reg[9][6]  ( .D(n341), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][6] ) );
  DFFARX1 \regf_reg[9][5]  ( .D(n340), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][5] ) );
  DFFARX1 \regf_reg[9][4]  ( .D(n339), .CLK(clk), .RSTB(n2681), .Q(
        \regf[9][4] ) );
  DFFARX1 \regf_reg[9][3]  ( .D(n338), .CLK(clk), .RSTB(n2682), .Q(
        \regf[9][3] ) );
  DFFARX1 \regf_reg[9][2]  ( .D(n337), .CLK(clk), .RSTB(n2682), .Q(
        \regf[9][2] ) );
  DFFARX1 \regf_reg[9][1]  ( .D(n336), .CLK(clk), .RSTB(n2682), .Q(
        \regf[9][1] ) );
  DFFARX1 \regf_reg[9][0]  ( .D(n335), .CLK(clk), .RSTB(n2682), .Q(
        \regf[9][0] ) );
  DFFARX1 \regf_reg[8][31]  ( .D(n334), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][31] ) );
  DFFARX1 \regf_reg[8][30]  ( .D(n333), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][30] ) );
  DFFARX1 \regf_reg[8][29]  ( .D(n332), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][29] ) );
  DFFARX1 \regf_reg[8][28]  ( .D(n331), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][28] ) );
  DFFARX1 \regf_reg[8][27]  ( .D(n330), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][27] ) );
  DFFARX1 \regf_reg[8][26]  ( .D(n329), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][26] ) );
  DFFARX1 \regf_reg[8][25]  ( .D(n328), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][25] ) );
  DFFARX1 \regf_reg[8][24]  ( .D(n327), .CLK(clk), .RSTB(n2682), .Q(
        \regf[8][24] ) );
  DFFARX1 \regf_reg[8][23]  ( .D(n326), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][23] ) );
  DFFARX1 \regf_reg[8][22]  ( .D(n325), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][22] ) );
  DFFARX1 \regf_reg[8][21]  ( .D(n324), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][21] ) );
  DFFARX1 \regf_reg[8][20]  ( .D(n323), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][20] ) );
  DFFARX1 \regf_reg[8][19]  ( .D(n322), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][19] ) );
  DFFARX1 \regf_reg[8][18]  ( .D(n321), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][18] ) );
  DFFARX1 \regf_reg[8][17]  ( .D(n320), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][17] ) );
  DFFARX1 \regf_reg[8][16]  ( .D(n319), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][16] ) );
  DFFARX1 \regf_reg[8][15]  ( .D(n318), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][15] ) );
  DFFARX1 \regf_reg[8][14]  ( .D(n317), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][14] ) );
  DFFARX1 \regf_reg[8][13]  ( .D(n316), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][13] ) );
  DFFARX1 \regf_reg[8][12]  ( .D(n315), .CLK(clk), .RSTB(n2683), .Q(
        \regf[8][12] ) );
  DFFARX1 \regf_reg[8][11]  ( .D(n314), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][11] ) );
  DFFARX1 \regf_reg[8][10]  ( .D(n313), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][10] ) );
  DFFARX1 \regf_reg[8][9]  ( .D(n312), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][9] ) );
  DFFARX1 \regf_reg[8][8]  ( .D(n311), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][8] ) );
  DFFARX1 \regf_reg[8][7]  ( .D(n310), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][7] ) );
  DFFARX1 \regf_reg[8][6]  ( .D(n309), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][6] ) );
  DFFARX1 \regf_reg[8][5]  ( .D(n308), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][5] ) );
  DFFARX1 \regf_reg[8][4]  ( .D(n307), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][4] ) );
  DFFARX1 \regf_reg[8][3]  ( .D(n306), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][3] ) );
  DFFARX1 \regf_reg[8][2]  ( .D(n305), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][2] ) );
  DFFARX1 \regf_reg[8][1]  ( .D(n304), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][1] ) );
  DFFARX1 \regf_reg[8][0]  ( .D(n303), .CLK(clk), .RSTB(n2684), .Q(
        \regf[8][0] ) );
  DFFARX1 \regf_reg[7][31]  ( .D(n302), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][31] ) );
  DFFARX1 \regf_reg[7][30]  ( .D(n301), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][30] ) );
  DFFARX1 \regf_reg[7][29]  ( .D(n300), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][29] ) );
  DFFARX1 \regf_reg[7][28]  ( .D(n299), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][28] ) );
  DFFARX1 \regf_reg[7][27]  ( .D(n298), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][27] ) );
  DFFARX1 \regf_reg[7][26]  ( .D(n297), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][26] ) );
  DFFARX1 \regf_reg[7][25]  ( .D(n296), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][25] ) );
  DFFARX1 \regf_reg[7][24]  ( .D(n295), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][24] ) );
  DFFARX1 \regf_reg[7][23]  ( .D(n294), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][23] ) );
  DFFARX1 \regf_reg[7][22]  ( .D(n293), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][22] ) );
  DFFARX1 \regf_reg[7][21]  ( .D(n292), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][21] ) );
  DFFARX1 \regf_reg[7][20]  ( .D(n291), .CLK(clk), .RSTB(n2685), .Q(
        \regf[7][20] ) );
  DFFARX1 \regf_reg[7][19]  ( .D(n290), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][19] ) );
  DFFARX1 \regf_reg[7][18]  ( .D(n289), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][18] ) );
  DFFARX1 \regf_reg[7][17]  ( .D(n288), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][17] ) );
  DFFARX1 \regf_reg[7][16]  ( .D(n287), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][16] ) );
  DFFARX1 \regf_reg[7][15]  ( .D(n286), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][15] ) );
  DFFARX1 \regf_reg[7][14]  ( .D(n285), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][14] ) );
  DFFARX1 \regf_reg[7][13]  ( .D(n284), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][13] ) );
  DFFARX1 \regf_reg[7][12]  ( .D(n283), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][12] ) );
  DFFARX1 \regf_reg[7][11]  ( .D(n282), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][11] ) );
  DFFARX1 \regf_reg[7][10]  ( .D(n281), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][10] ) );
  DFFARX1 \regf_reg[7][9]  ( .D(n280), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][9] ) );
  DFFARX1 \regf_reg[7][8]  ( .D(n279), .CLK(clk), .RSTB(n2686), .Q(
        \regf[7][8] ) );
  DFFARX1 \regf_reg[7][7]  ( .D(n278), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][7] ) );
  DFFARX1 \regf_reg[7][6]  ( .D(n277), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][6] ) );
  DFFARX1 \regf_reg[7][5]  ( .D(n276), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][5] ) );
  DFFARX1 \regf_reg[7][4]  ( .D(n275), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][4] ) );
  DFFARX1 \regf_reg[7][3]  ( .D(n274), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][3] ) );
  DFFARX1 \regf_reg[7][2]  ( .D(n273), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][2] ) );
  DFFARX1 \regf_reg[7][1]  ( .D(n272), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][1] ) );
  DFFARX1 \regf_reg[7][0]  ( .D(n271), .CLK(clk), .RSTB(n2687), .Q(
        \regf[7][0] ) );
  DFFARX1 \regf_reg[6][31]  ( .D(n270), .CLK(clk), .RSTB(n2687), .Q(
        \regf[6][31] ) );
  DFFARX1 \regf_reg[6][30]  ( .D(n269), .CLK(clk), .RSTB(n2687), .Q(
        \regf[6][30] ) );
  DFFARX1 \regf_reg[6][29]  ( .D(n268), .CLK(clk), .RSTB(n2687), .Q(
        \regf[6][29] ) );
  DFFARX1 \regf_reg[6][28]  ( .D(n267), .CLK(clk), .RSTB(n2687), .Q(
        \regf[6][28] ) );
  DFFARX1 \regf_reg[6][27]  ( .D(n266), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][27] ) );
  DFFARX1 \regf_reg[6][26]  ( .D(n265), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][26] ) );
  DFFARX1 \regf_reg[6][25]  ( .D(n264), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][25] ) );
  DFFARX1 \regf_reg[6][24]  ( .D(n263), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][24] ) );
  DFFARX1 \regf_reg[6][23]  ( .D(n262), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][23] ) );
  DFFARX1 \regf_reg[6][22]  ( .D(n261), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][22] ) );
  DFFARX1 \regf_reg[6][21]  ( .D(n260), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][21] ) );
  DFFARX1 \regf_reg[6][20]  ( .D(n259), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][20] ) );
  DFFARX1 \regf_reg[6][19]  ( .D(n258), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][19] ) );
  DFFARX1 \regf_reg[6][18]  ( .D(n257), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][18] ) );
  DFFARX1 \regf_reg[6][17]  ( .D(n256), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][17] ) );
  DFFARX1 \regf_reg[6][16]  ( .D(n255), .CLK(clk), .RSTB(n2688), .Q(
        \regf[6][16] ) );
  DFFARX1 \regf_reg[6][15]  ( .D(n254), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][15] ) );
  DFFARX1 \regf_reg[6][14]  ( .D(n253), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][14] ) );
  DFFARX1 \regf_reg[6][13]  ( .D(n252), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][13] ) );
  DFFARX1 \regf_reg[6][12]  ( .D(n251), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][12] ) );
  DFFARX1 \regf_reg[6][11]  ( .D(n250), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][11] ) );
  DFFARX1 \regf_reg[6][10]  ( .D(n249), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][10] ) );
  DFFARX1 \regf_reg[6][9]  ( .D(n248), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][9] ) );
  DFFARX1 \regf_reg[6][8]  ( .D(n247), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][8] ) );
  DFFARX1 \regf_reg[6][7]  ( .D(n246), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][7] ) );
  DFFARX1 \regf_reg[6][6]  ( .D(n245), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][6] ) );
  DFFARX1 \regf_reg[6][5]  ( .D(n244), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][5] ) );
  DFFARX1 \regf_reg[6][4]  ( .D(n243), .CLK(clk), .RSTB(n2689), .Q(
        \regf[6][4] ) );
  DFFARX1 \regf_reg[6][3]  ( .D(n242), .CLK(clk), .RSTB(n2690), .Q(
        \regf[6][3] ) );
  DFFARX1 \regf_reg[6][2]  ( .D(n241), .CLK(clk), .RSTB(n2690), .Q(
        \regf[6][2] ) );
  DFFARX1 \regf_reg[6][1]  ( .D(n240), .CLK(clk), .RSTB(n2690), .Q(
        \regf[6][1] ) );
  DFFARX1 \regf_reg[6][0]  ( .D(n239), .CLK(clk), .RSTB(n2690), .Q(
        \regf[6][0] ) );
  DFFARX1 \regf_reg[5][31]  ( .D(n238), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][31] ) );
  DFFARX1 \regf_reg[5][30]  ( .D(n237), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][30] ) );
  DFFARX1 \regf_reg[5][29]  ( .D(n236), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][29] ) );
  DFFARX1 \regf_reg[5][28]  ( .D(n235), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][28] ) );
  DFFARX1 \regf_reg[5][27]  ( .D(n234), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][27] ) );
  DFFARX1 \regf_reg[5][26]  ( .D(n233), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][26] ) );
  DFFARX1 \regf_reg[5][25]  ( .D(n232), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][25] ) );
  DFFARX1 \regf_reg[5][24]  ( .D(n231), .CLK(clk), .RSTB(n2690), .Q(
        \regf[5][24] ) );
  DFFARX1 \regf_reg[5][23]  ( .D(n230), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][23] ) );
  DFFARX1 \regf_reg[5][22]  ( .D(n229), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][22] ) );
  DFFARX1 \regf_reg[5][21]  ( .D(n228), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][21] ) );
  DFFARX1 \regf_reg[5][20]  ( .D(n227), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][20] ) );
  DFFARX1 \regf_reg[5][19]  ( .D(n226), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][19] ) );
  DFFARX1 \regf_reg[5][18]  ( .D(n225), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][18] ) );
  DFFARX1 \regf_reg[5][17]  ( .D(n224), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][17] ) );
  DFFARX1 \regf_reg[5][16]  ( .D(n223), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][16] ) );
  DFFARX1 \regf_reg[5][15]  ( .D(n222), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][15] ) );
  DFFARX1 \regf_reg[5][14]  ( .D(n221), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][14] ) );
  DFFARX1 \regf_reg[5][13]  ( .D(n220), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][13] ) );
  DFFARX1 \regf_reg[5][12]  ( .D(n219), .CLK(clk), .RSTB(n2691), .Q(
        \regf[5][12] ) );
  DFFARX1 \regf_reg[5][11]  ( .D(n218), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][11] ) );
  DFFARX1 \regf_reg[5][10]  ( .D(n217), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][10] ) );
  DFFARX1 \regf_reg[5][9]  ( .D(n216), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][9] ) );
  DFFARX1 \regf_reg[5][8]  ( .D(n215), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][8] ) );
  DFFARX1 \regf_reg[5][7]  ( .D(n214), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][7] ) );
  DFFARX1 \regf_reg[5][6]  ( .D(n213), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][6] ) );
  DFFARX1 \regf_reg[5][5]  ( .D(n212), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][5] ) );
  DFFARX1 \regf_reg[5][4]  ( .D(n211), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][4] ) );
  DFFARX1 \regf_reg[5][3]  ( .D(n210), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][3] ) );
  DFFARX1 \regf_reg[5][2]  ( .D(n209), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][2] ) );
  DFFARX1 \regf_reg[5][1]  ( .D(n208), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][1] ) );
  DFFARX1 \regf_reg[5][0]  ( .D(n207), .CLK(clk), .RSTB(n2692), .Q(
        \regf[5][0] ) );
  DFFARX1 \regf_reg[4][31]  ( .D(n206), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][31] ) );
  DFFARX1 \regf_reg[4][30]  ( .D(n205), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][30] ) );
  DFFARX1 \regf_reg[4][29]  ( .D(n204), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][29] ) );
  DFFARX1 \regf_reg[4][28]  ( .D(n203), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][28] ) );
  DFFARX1 \regf_reg[4][27]  ( .D(n202), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][27] ) );
  DFFARX1 \regf_reg[4][26]  ( .D(n201), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][26] ) );
  DFFARX1 \regf_reg[4][25]  ( .D(n200), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][25] ) );
  DFFARX1 \regf_reg[4][24]  ( .D(n199), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][24] ) );
  DFFARX1 \regf_reg[4][23]  ( .D(n198), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][23] ) );
  DFFARX1 \regf_reg[4][22]  ( .D(n197), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][22] ) );
  DFFARX1 \regf_reg[4][21]  ( .D(n196), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][21] ) );
  DFFARX1 \regf_reg[4][20]  ( .D(n195), .CLK(clk), .RSTB(n2693), .Q(
        \regf[4][20] ) );
  DFFARX1 \regf_reg[4][19]  ( .D(n194), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][19] ) );
  DFFARX1 \regf_reg[4][18]  ( .D(n193), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][18] ) );
  DFFARX1 \regf_reg[4][17]  ( .D(n192), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][17] ) );
  DFFARX1 \regf_reg[4][16]  ( .D(n191), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][16] ) );
  DFFARX1 \regf_reg[4][15]  ( .D(n190), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][15] ) );
  DFFARX1 \regf_reg[4][14]  ( .D(n189), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][14] ) );
  DFFARX1 \regf_reg[4][13]  ( .D(n188), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][13] ) );
  DFFARX1 \regf_reg[4][12]  ( .D(n187), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][12] ) );
  DFFARX1 \regf_reg[4][11]  ( .D(n186), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][11] ) );
  DFFARX1 \regf_reg[4][10]  ( .D(n185), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][10] ) );
  DFFARX1 \regf_reg[4][9]  ( .D(n184), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][9] ) );
  DFFARX1 \regf_reg[4][8]  ( .D(n183), .CLK(clk), .RSTB(n2694), .Q(
        \regf[4][8] ) );
  DFFARX1 \regf_reg[4][7]  ( .D(n182), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][7] ) );
  DFFARX1 \regf_reg[4][6]  ( .D(n181), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][6] ) );
  DFFARX1 \regf_reg[4][5]  ( .D(n180), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][5] ) );
  DFFARX1 \regf_reg[4][4]  ( .D(n179), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][4] ) );
  DFFARX1 \regf_reg[4][3]  ( .D(n178), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][3] ) );
  DFFARX1 \regf_reg[4][2]  ( .D(n177), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][2] ) );
  DFFARX1 \regf_reg[4][1]  ( .D(n176), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][1] ) );
  DFFARX1 \regf_reg[4][0]  ( .D(n175), .CLK(clk), .RSTB(n2695), .Q(
        \regf[4][0] ) );
  DFFARX1 \regf_reg[3][31]  ( .D(n174), .CLK(clk), .RSTB(n2695), .Q(
        \regf[3][31] ) );
  DFFARX1 \regf_reg[3][30]  ( .D(n173), .CLK(clk), .RSTB(n2695), .Q(
        \regf[3][30] ) );
  DFFARX1 \regf_reg[3][29]  ( .D(n172), .CLK(clk), .RSTB(n2695), .Q(
        \regf[3][29] ) );
  DFFARX1 \regf_reg[3][28]  ( .D(n171), .CLK(clk), .RSTB(n2695), .Q(
        \regf[3][28] ) );
  DFFARX1 \regf_reg[3][27]  ( .D(n170), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][27] ) );
  DFFARX1 \regf_reg[3][26]  ( .D(n169), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][26] ) );
  DFFARX1 \regf_reg[3][25]  ( .D(n168), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][25] ) );
  DFFARX1 \regf_reg[3][24]  ( .D(n167), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][24] ) );
  DFFARX1 \regf_reg[3][23]  ( .D(n166), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][23] ) );
  DFFARX1 \regf_reg[3][22]  ( .D(n165), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][22] ) );
  DFFARX1 \regf_reg[3][21]  ( .D(n164), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][21] ) );
  DFFARX1 \regf_reg[3][20]  ( .D(n163), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][20] ) );
  DFFARX1 \regf_reg[3][19]  ( .D(n162), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][19] ) );
  DFFARX1 \regf_reg[3][18]  ( .D(n161), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][18] ) );
  DFFARX1 \regf_reg[3][17]  ( .D(n160), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][17] ) );
  DFFARX1 \regf_reg[3][16]  ( .D(n159), .CLK(clk), .RSTB(n2696), .Q(
        \regf[3][16] ) );
  DFFARX1 \regf_reg[3][15]  ( .D(n158), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][15] ) );
  DFFARX1 \regf_reg[3][14]  ( .D(n157), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][14] ) );
  DFFARX1 \regf_reg[3][13]  ( .D(n156), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][13] ) );
  DFFARX1 \regf_reg[3][12]  ( .D(n155), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][12] ) );
  DFFARX1 \regf_reg[3][11]  ( .D(n154), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][11] ) );
  DFFARX1 \regf_reg[3][10]  ( .D(n153), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][10] ) );
  DFFARX1 \regf_reg[3][9]  ( .D(n152), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][9] ) );
  DFFARX1 \regf_reg[3][8]  ( .D(n151), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][8] ) );
  DFFARX1 \regf_reg[3][7]  ( .D(n150), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][7] ) );
  DFFARX1 \regf_reg[3][6]  ( .D(n149), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][6] ) );
  DFFARX1 \regf_reg[3][5]  ( .D(n148), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][5] ) );
  DFFARX1 \regf_reg[3][4]  ( .D(n147), .CLK(clk), .RSTB(n2697), .Q(
        \regf[3][4] ) );
  DFFARX1 \regf_reg[3][3]  ( .D(n146), .CLK(clk), .RSTB(n2698), .Q(
        \regf[3][3] ) );
  DFFARX1 \regf_reg[3][2]  ( .D(n145), .CLK(clk), .RSTB(n2698), .Q(
        \regf[3][2] ) );
  DFFARX1 \regf_reg[3][1]  ( .D(n144), .CLK(clk), .RSTB(n2698), .Q(
        \regf[3][1] ) );
  DFFARX1 \regf_reg[3][0]  ( .D(n143), .CLK(clk), .RSTB(n2698), .Q(
        \regf[3][0] ) );
  DFFARX1 \regf_reg[2][31]  ( .D(n142), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][31] ) );
  DFFARX1 \regf_reg[2][30]  ( .D(n141), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][30] ) );
  DFFARX1 \regf_reg[2][29]  ( .D(n140), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][29] ) );
  DFFARX1 \regf_reg[2][28]  ( .D(n139), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][28] ) );
  DFFARX1 \regf_reg[2][27]  ( .D(n138), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][27] ) );
  DFFARX1 \regf_reg[2][26]  ( .D(n137), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][26] ) );
  DFFARX1 \regf_reg[2][25]  ( .D(n136), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][25] ), .QN(n1098) );
  DFFARX1 \regf_reg[2][24]  ( .D(n135), .CLK(clk), .RSTB(n2698), .Q(
        \regf[2][24] ) );
  DFFARX1 \regf_reg[2][23]  ( .D(n134), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][23] ) );
  DFFARX1 \regf_reg[2][22]  ( .D(n133), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][22] ), .QN(n1144) );
  DFFARX1 \regf_reg[2][21]  ( .D(n132), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][21] ) );
  DFFARX1 \regf_reg[2][20]  ( .D(n131), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][20] ) );
  DFFARX1 \regf_reg[2][19]  ( .D(n130), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][19] ) );
  DFFARX1 \regf_reg[2][18]  ( .D(n129), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][18] ) );
  DFFARX1 \regf_reg[2][17]  ( .D(n128), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][17] ) );
  DFFARX1 \regf_reg[2][16]  ( .D(n127), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][16] ) );
  DFFARX1 \regf_reg[2][15]  ( .D(n126), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][15] ) );
  DFFARX1 \regf_reg[2][14]  ( .D(n125), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][14] ), .QN(n1136) );
  DFFARX1 \regf_reg[2][13]  ( .D(n124), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][13] ) );
  DFFARX1 \regf_reg[2][12]  ( .D(n123), .CLK(clk), .RSTB(n2699), .Q(
        \regf[2][12] ), .QN(n1122) );
  DFFARX1 \regf_reg[2][11]  ( .D(n122), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][11] ) );
  DFFARX1 \regf_reg[2][10]  ( .D(n121), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][10] ) );
  DFFARX1 \regf_reg[2][9]  ( .D(n120), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][9] ) );
  DFFARX1 \regf_reg[2][8]  ( .D(n119), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][8] ) );
  DFFARX1 \regf_reg[2][7]  ( .D(n118), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][7] ) );
  DFFARX1 \regf_reg[2][6]  ( .D(n117), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][6] ), .QN(n1118) );
  DFFARX1 \regf_reg[2][5]  ( .D(n116), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][5] ), .QN(n1100) );
  DFFARX1 \regf_reg[2][4]  ( .D(n115), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][4] ) );
  DFFARX1 \regf_reg[2][3]  ( .D(n114), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][3] ), .QN(n1099) );
  DFFARX1 \regf_reg[2][2]  ( .D(n113), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][2] ) );
  DFFARX1 \regf_reg[2][1]  ( .D(n112), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][1] ), .QN(n1102) );
  DFFARX1 \regf_reg[2][0]  ( .D(n111), .CLK(clk), .RSTB(n2700), .Q(
        \regf[2][0] ) );
  DFFARX1 \regf_reg[1][31]  ( .D(n110), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][31] ) );
  DFFARX1 \regf_reg[1][30]  ( .D(n109), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][30] ) );
  DFFARX1 \regf_reg[1][29]  ( .D(n108), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][29] ) );
  DFFARX1 \regf_reg[1][28]  ( .D(n107), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][28] ) );
  DFFARX1 \regf_reg[1][27]  ( .D(n106), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][27] ) );
  DFFARX1 \regf_reg[1][26]  ( .D(n105), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][26] ) );
  DFFARX1 \regf_reg[1][25]  ( .D(n104), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][25] ) );
  DFFARX1 \regf_reg[1][24]  ( .D(n103), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][24] ) );
  DFFARX1 \regf_reg[1][23]  ( .D(n102), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][23] ) );
  DFFARX1 \regf_reg[1][22]  ( .D(n101), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][22] ) );
  DFFARX1 \regf_reg[1][21]  ( .D(n100), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][21] ) );
  DFFARX1 \regf_reg[1][20]  ( .D(n99), .CLK(clk), .RSTB(n2701), .Q(
        \regf[1][20] ) );
  DFFARX1 \regf_reg[1][19]  ( .D(n98), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][19] ) );
  DFFARX1 \regf_reg[1][18]  ( .D(n97), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][18] ) );
  DFFARX1 \regf_reg[1][17]  ( .D(n96), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][17] ) );
  DFFARX1 \regf_reg[1][16]  ( .D(n95), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][16] ) );
  DFFARX1 \regf_reg[1][15]  ( .D(n94), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][15] ) );
  DFFARX1 \regf_reg[1][14]  ( .D(n93), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][14] ) );
  DFFARX1 \regf_reg[1][13]  ( .D(n92), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][13] ) );
  DFFARX1 \regf_reg[1][12]  ( .D(n91), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][12] ) );
  DFFARX1 \regf_reg[1][11]  ( .D(n90), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][11] ) );
  DFFARX1 \regf_reg[1][10]  ( .D(n89), .CLK(clk), .RSTB(n2702), .Q(
        \regf[1][10] ) );
  DFFARX1 \regf_reg[1][9]  ( .D(n88), .CLK(clk), .RSTB(n2702), .Q(\regf[1][9] ) );
  DFFARX1 \regf_reg[1][8]  ( .D(n87), .CLK(clk), .RSTB(n2702), .Q(\regf[1][8] ) );
  DFFARX1 \regf_reg[1][7]  ( .D(n86), .CLK(clk), .RSTB(n2703), .Q(\regf[1][7] ) );
  DFFARX1 \regf_reg[1][6]  ( .D(n85), .CLK(clk), .RSTB(n2703), .Q(\regf[1][6] ) );
  DFFARX1 \regf_reg[1][5]  ( .D(n84), .CLK(clk), .RSTB(n2703), .Q(\regf[1][5] ) );
  DFFARX1 \regf_reg[1][4]  ( .D(n83), .CLK(clk), .RSTB(n2703), .Q(\regf[1][4] ) );
  DFFARX1 \regf_reg[1][3]  ( .D(n82), .CLK(clk), .RSTB(n2703), .Q(\regf[1][3] ) );
  DFFARX1 \regf_reg[1][2]  ( .D(n81), .CLK(clk), .RSTB(n2703), .Q(\regf[1][2] ) );
  DFFARX1 \regf_reg[1][1]  ( .D(n80), .CLK(clk), .RSTB(n2703), .Q(\regf[1][1] ) );
  DFFARX1 \regf_reg[1][0]  ( .D(n79), .CLK(clk), .RSTB(n2703), .Q(\regf[1][0] ) );
  AO22X1 U100 ( .IN1(n2525), .IN2(n2522), .IN3(\regf[1][0] ), .IN4(n2521), .Q(
        n79) );
  AO22X1 U101 ( .IN1(n2528), .IN2(n2522), .IN3(\regf[1][1] ), .IN4(n2521), .Q(
        n80) );
  AO22X1 U102 ( .IN1(n2531), .IN2(n2522), .IN3(\regf[1][2] ), .IN4(n2521), .Q(
        n81) );
  AO22X1 U103 ( .IN1(n2534), .IN2(n2522), .IN3(\regf[1][3] ), .IN4(n2521), .Q(
        n82) );
  AO22X1 U104 ( .IN1(n2537), .IN2(n2523), .IN3(\regf[1][4] ), .IN4(n2521), .Q(
        n83) );
  AO22X1 U105 ( .IN1(n2540), .IN2(n2524), .IN3(\regf[1][5] ), .IN4(n2521), .Q(
        n84) );
  AO22X1 U106 ( .IN1(n2543), .IN2(n2523), .IN3(\regf[1][6] ), .IN4(n2521), .Q(
        n85) );
  AO22X1 U107 ( .IN1(n2546), .IN2(n2523), .IN3(\regf[1][7] ), .IN4(n2521), .Q(
        n86) );
  AO22X1 U108 ( .IN1(n2549), .IN2(n2524), .IN3(\regf[1][8] ), .IN4(n2521), .Q(
        n87) );
  AO22X1 U109 ( .IN1(n2552), .IN2(n2524), .IN3(\regf[1][9] ), .IN4(n2521), .Q(
        n88) );
  AO22X1 U110 ( .IN1(n2555), .IN2(n2523), .IN3(\regf[1][10] ), .IN4(n2521), 
        .Q(n89) );
  AO22X1 U111 ( .IN1(n2558), .IN2(n2523), .IN3(\regf[1][11] ), .IN4(n2521), 
        .Q(n90) );
  AO22X1 U112 ( .IN1(n2561), .IN2(n2523), .IN3(\regf[1][12] ), .IN4(n2521), 
        .Q(n91) );
  AO22X1 U113 ( .IN1(n2564), .IN2(n2523), .IN3(\regf[1][13] ), .IN4(n2520), 
        .Q(n92) );
  AO22X1 U114 ( .IN1(n2567), .IN2(n2523), .IN3(\regf[1][14] ), .IN4(n37), .Q(
        n93) );
  AO22X1 U115 ( .IN1(n2570), .IN2(n2523), .IN3(\regf[1][15] ), .IN4(n37), .Q(
        n94) );
  AO22X1 U116 ( .IN1(n2573), .IN2(n2523), .IN3(\regf[1][16] ), .IN4(n37), .Q(
        n95) );
  AO22X1 U117 ( .IN1(n2576), .IN2(n2523), .IN3(\regf[1][17] ), .IN4(n37), .Q(
        n96) );
  AO22X1 U118 ( .IN1(n2579), .IN2(n2524), .IN3(\regf[1][18] ), .IN4(n37), .Q(
        n97) );
  AO22X1 U119 ( .IN1(n2582), .IN2(n2523), .IN3(\regf[1][19] ), .IN4(n37), .Q(
        n98) );
  AO22X1 U120 ( .IN1(n2585), .IN2(n2524), .IN3(\regf[1][20] ), .IN4(n2520), 
        .Q(n99) );
  AO22X1 U121 ( .IN1(n2588), .IN2(n2523), .IN3(\regf[1][21] ), .IN4(n2520), 
        .Q(n100) );
  AO22X1 U122 ( .IN1(n2591), .IN2(n2524), .IN3(\regf[1][22] ), .IN4(n2520), 
        .Q(n101) );
  AO22X1 U123 ( .IN1(n2594), .IN2(n2523), .IN3(\regf[1][23] ), .IN4(n2520), 
        .Q(n102) );
  AO22X1 U124 ( .IN1(n2597), .IN2(n2524), .IN3(\regf[1][24] ), .IN4(n2520), 
        .Q(n103) );
  AO22X1 U125 ( .IN1(n2600), .IN2(n2524), .IN3(\regf[1][25] ), .IN4(n2520), 
        .Q(n104) );
  AO22X1 U126 ( .IN1(n2603), .IN2(n2524), .IN3(\regf[1][26] ), .IN4(n2520), 
        .Q(n105) );
  AO22X1 U127 ( .IN1(n2606), .IN2(n2524), .IN3(\regf[1][27] ), .IN4(n2520), 
        .Q(n106) );
  AO22X1 U128 ( .IN1(n2609), .IN2(n2524), .IN3(\regf[1][28] ), .IN4(n2520), 
        .Q(n107) );
  AO22X1 U129 ( .IN1(n2612), .IN2(n2524), .IN3(\regf[1][29] ), .IN4(n2520), 
        .Q(n108) );
  AO22X1 U130 ( .IN1(n2615), .IN2(n2524), .IN3(\regf[1][30] ), .IN4(n2520), 
        .Q(n109) );
  AO22X1 U131 ( .IN1(n2618), .IN2(n2524), .IN3(\regf[1][31] ), .IN4(n2520), 
        .Q(n110) );
  AO22X1 U132 ( .IN1(n2517), .IN2(n2525), .IN3(\regf[2][0] ), .IN4(n2516), .Q(
        n111) );
  AO22X1 U133 ( .IN1(n2517), .IN2(n2528), .IN3(\regf[2][1] ), .IN4(n2516), .Q(
        n112) );
  AO22X1 U134 ( .IN1(n2517), .IN2(n2531), .IN3(\regf[2][2] ), .IN4(n2516), .Q(
        n113) );
  AO22X1 U135 ( .IN1(n2517), .IN2(n2534), .IN3(\regf[2][3] ), .IN4(n2516), .Q(
        n114) );
  AO22X1 U136 ( .IN1(n2518), .IN2(n2537), .IN3(\regf[2][4] ), .IN4(n2516), .Q(
        n115) );
  AO22X1 U137 ( .IN1(n2519), .IN2(n2540), .IN3(\regf[2][5] ), .IN4(n2516), .Q(
        n116) );
  AO22X1 U138 ( .IN1(n2518), .IN2(n2543), .IN3(\regf[2][6] ), .IN4(n2516), .Q(
        n117) );
  AO22X1 U139 ( .IN1(n2518), .IN2(n2546), .IN3(\regf[2][7] ), .IN4(n2516), .Q(
        n118) );
  AO22X1 U140 ( .IN1(n2519), .IN2(n2549), .IN3(\regf[2][8] ), .IN4(n2516), .Q(
        n119) );
  AO22X1 U141 ( .IN1(n2519), .IN2(n2552), .IN3(\regf[2][9] ), .IN4(n2516), .Q(
        n120) );
  AO22X1 U142 ( .IN1(n2518), .IN2(n2555), .IN3(\regf[2][10] ), .IN4(n2516), 
        .Q(n121) );
  AO22X1 U143 ( .IN1(n2518), .IN2(n2558), .IN3(\regf[2][11] ), .IN4(n2515), 
        .Q(n122) );
  AO22X1 U144 ( .IN1(n2518), .IN2(n2561), .IN3(\regf[2][12] ), .IN4(n40), .Q(
        n123) );
  AO22X1 U145 ( .IN1(n2518), .IN2(n2564), .IN3(\regf[2][13] ), .IN4(n40), .Q(
        n124) );
  AO22X1 U146 ( .IN1(n2518), .IN2(n2567), .IN3(\regf[2][14] ), .IN4(n40), .Q(
        n125) );
  AO22X1 U147 ( .IN1(n2518), .IN2(n2570), .IN3(\regf[2][15] ), .IN4(n40), .Q(
        n126) );
  AO22X1 U148 ( .IN1(n2518), .IN2(n2573), .IN3(\regf[2][16] ), .IN4(n40), .Q(
        n127) );
  AO22X1 U149 ( .IN1(n2518), .IN2(n2576), .IN3(\regf[2][17] ), .IN4(n40), .Q(
        n128) );
  AO22X1 U150 ( .IN1(n2519), .IN2(n2579), .IN3(\regf[2][18] ), .IN4(n2516), 
        .Q(n129) );
  AO22X1 U151 ( .IN1(n2518), .IN2(n2582), .IN3(\regf[2][19] ), .IN4(n2516), 
        .Q(n130) );
  AO22X1 U152 ( .IN1(n2519), .IN2(n2585), .IN3(\regf[2][20] ), .IN4(n2515), 
        .Q(n131) );
  AO22X1 U153 ( .IN1(n2518), .IN2(n2588), .IN3(\regf[2][21] ), .IN4(n2515), 
        .Q(n132) );
  AO22X1 U154 ( .IN1(n2519), .IN2(n2591), .IN3(\regf[2][22] ), .IN4(n2515), 
        .Q(n133) );
  AO22X1 U155 ( .IN1(n2518), .IN2(n2594), .IN3(\regf[2][23] ), .IN4(n2515), 
        .Q(n134) );
  AO22X1 U156 ( .IN1(n2519), .IN2(n2597), .IN3(\regf[2][24] ), .IN4(n2515), 
        .Q(n135) );
  AO22X1 U157 ( .IN1(n2519), .IN2(n2600), .IN3(\regf[2][25] ), .IN4(n2515), 
        .Q(n136) );
  AO22X1 U158 ( .IN1(n2519), .IN2(n2603), .IN3(\regf[2][26] ), .IN4(n2515), 
        .Q(n137) );
  AO22X1 U159 ( .IN1(n2519), .IN2(n2606), .IN3(\regf[2][27] ), .IN4(n2515), 
        .Q(n138) );
  AO22X1 U160 ( .IN1(n2519), .IN2(n2609), .IN3(\regf[2][28] ), .IN4(n2515), 
        .Q(n139) );
  AO22X1 U161 ( .IN1(n2519), .IN2(n2612), .IN3(\regf[2][29] ), .IN4(n2515), 
        .Q(n140) );
  AO22X1 U162 ( .IN1(n2519), .IN2(n2615), .IN3(\regf[2][30] ), .IN4(n2515), 
        .Q(n141) );
  AO22X1 U163 ( .IN1(n2519), .IN2(n2618), .IN3(\regf[2][31] ), .IN4(n2515), 
        .Q(n142) );
  AO22X1 U164 ( .IN1(n2512), .IN2(n2525), .IN3(\regf[3][0] ), .IN4(n2511), .Q(
        n143) );
  AO22X1 U165 ( .IN1(n2512), .IN2(n2528), .IN3(\regf[3][1] ), .IN4(n2511), .Q(
        n144) );
  AO22X1 U166 ( .IN1(n2512), .IN2(n2531), .IN3(\regf[3][2] ), .IN4(n2511), .Q(
        n145) );
  AO22X1 U167 ( .IN1(n2512), .IN2(n2534), .IN3(\regf[3][3] ), .IN4(n2511), .Q(
        n146) );
  AO22X1 U168 ( .IN1(n2514), .IN2(n2537), .IN3(\regf[3][4] ), .IN4(n2511), .Q(
        n147) );
  AO22X1 U169 ( .IN1(n2513), .IN2(n2540), .IN3(\regf[3][5] ), .IN4(n2511), .Q(
        n148) );
  AO22X1 U170 ( .IN1(n2513), .IN2(n2543), .IN3(\regf[3][6] ), .IN4(n2511), .Q(
        n149) );
  AO22X1 U171 ( .IN1(n2514), .IN2(n2546), .IN3(\regf[3][7] ), .IN4(n2511), .Q(
        n150) );
  AO22X1 U172 ( .IN1(n2513), .IN2(n2549), .IN3(\regf[3][8] ), .IN4(n2511), .Q(
        n151) );
  AO22X1 U173 ( .IN1(n2513), .IN2(n2552), .IN3(\regf[3][9] ), .IN4(n2511), .Q(
        n152) );
  AO22X1 U174 ( .IN1(n2514), .IN2(n2555), .IN3(\regf[3][10] ), .IN4(n2511), 
        .Q(n153) );
  AO22X1 U175 ( .IN1(n2514), .IN2(n2558), .IN3(\regf[3][11] ), .IN4(n2511), 
        .Q(n154) );
  AO22X1 U176 ( .IN1(n2513), .IN2(n2561), .IN3(\regf[3][12] ), .IN4(n2511), 
        .Q(n155) );
  AO22X1 U177 ( .IN1(n2514), .IN2(n2564), .IN3(\regf[3][13] ), .IN4(n2510), 
        .Q(n156) );
  AO22X1 U178 ( .IN1(n2513), .IN2(n2567), .IN3(\regf[3][14] ), .IN4(n42), .Q(
        n157) );
  AO22X1 U179 ( .IN1(n2514), .IN2(n2570), .IN3(\regf[3][15] ), .IN4(n42), .Q(
        n158) );
  AO22X1 U180 ( .IN1(n2513), .IN2(n2573), .IN3(\regf[3][16] ), .IN4(n42), .Q(
        n159) );
  AO22X1 U181 ( .IN1(n2514), .IN2(n2576), .IN3(\regf[3][17] ), .IN4(n42), .Q(
        n160) );
  AO22X1 U182 ( .IN1(n2513), .IN2(n2579), .IN3(\regf[3][18] ), .IN4(n42), .Q(
        n161) );
  AO22X1 U183 ( .IN1(n2513), .IN2(n2582), .IN3(\regf[3][19] ), .IN4(n42), .Q(
        n162) );
  AO22X1 U184 ( .IN1(n2513), .IN2(n2585), .IN3(\regf[3][20] ), .IN4(n2510), 
        .Q(n163) );
  AO22X1 U185 ( .IN1(n2513), .IN2(n2588), .IN3(\regf[3][21] ), .IN4(n2510), 
        .Q(n164) );
  AO22X1 U186 ( .IN1(n2513), .IN2(n2591), .IN3(\regf[3][22] ), .IN4(n2510), 
        .Q(n165) );
  AO22X1 U187 ( .IN1(n2513), .IN2(n2594), .IN3(\regf[3][23] ), .IN4(n2510), 
        .Q(n166) );
  AO22X1 U188 ( .IN1(n2513), .IN2(n2597), .IN3(\regf[3][24] ), .IN4(n2510), 
        .Q(n167) );
  AO22X1 U189 ( .IN1(n2514), .IN2(n2600), .IN3(\regf[3][25] ), .IN4(n2510), 
        .Q(n168) );
  AO22X1 U190 ( .IN1(n2514), .IN2(n2603), .IN3(\regf[3][26] ), .IN4(n2510), 
        .Q(n169) );
  AO22X1 U191 ( .IN1(n2514), .IN2(n2606), .IN3(\regf[3][27] ), .IN4(n2510), 
        .Q(n170) );
  AO22X1 U192 ( .IN1(n2514), .IN2(n2609), .IN3(\regf[3][28] ), .IN4(n2510), 
        .Q(n171) );
  AO22X1 U193 ( .IN1(n2514), .IN2(n2612), .IN3(\regf[3][29] ), .IN4(n2510), 
        .Q(n172) );
  AO22X1 U194 ( .IN1(n2514), .IN2(n2615), .IN3(\regf[3][30] ), .IN4(n2510), 
        .Q(n173) );
  AO22X1 U195 ( .IN1(n2514), .IN2(n2618), .IN3(\regf[3][31] ), .IN4(n2510), 
        .Q(n174) );
  AO22X1 U196 ( .IN1(n2509), .IN2(n2525), .IN3(\regf[4][0] ), .IN4(n2507), .Q(
        n175) );
  AO22X1 U197 ( .IN1(n2508), .IN2(n2528), .IN3(\regf[4][1] ), .IN4(n2507), .Q(
        n176) );
  AO22X1 U198 ( .IN1(n2509), .IN2(n2531), .IN3(\regf[4][2] ), .IN4(n2507), .Q(
        n177) );
  AO22X1 U199 ( .IN1(n2508), .IN2(n2534), .IN3(\regf[4][3] ), .IN4(n2507), .Q(
        n178) );
  AO22X1 U200 ( .IN1(n2508), .IN2(n2537), .IN3(\regf[4][4] ), .IN4(n2507), .Q(
        n179) );
  AO22X1 U201 ( .IN1(n2509), .IN2(n2540), .IN3(\regf[4][5] ), .IN4(n2507), .Q(
        n180) );
  AO22X1 U202 ( .IN1(n2508), .IN2(n2543), .IN3(\regf[4][6] ), .IN4(n2507), .Q(
        n181) );
  AO22X1 U203 ( .IN1(n2508), .IN2(n2546), .IN3(\regf[4][7] ), .IN4(n2507), .Q(
        n182) );
  AO22X1 U204 ( .IN1(n2509), .IN2(n2549), .IN3(\regf[4][8] ), .IN4(n2507), .Q(
        n183) );
  AO22X1 U205 ( .IN1(n2509), .IN2(n2552), .IN3(\regf[4][9] ), .IN4(n2507), .Q(
        n184) );
  AO22X1 U206 ( .IN1(n2508), .IN2(n2555), .IN3(\regf[4][10] ), .IN4(n2507), 
        .Q(n185) );
  AO22X1 U207 ( .IN1(n2508), .IN2(n2558), .IN3(\regf[4][11] ), .IN4(n2507), 
        .Q(n186) );
  AO22X1 U208 ( .IN1(n2508), .IN2(n2561), .IN3(\regf[4][12] ), .IN4(n2507), 
        .Q(n187) );
  AO22X1 U209 ( .IN1(n2508), .IN2(n2564), .IN3(\regf[4][13] ), .IN4(n2506), 
        .Q(n188) );
  AO22X1 U210 ( .IN1(n2508), .IN2(n2567), .IN3(\regf[4][14] ), .IN4(n44), .Q(
        n189) );
  AO22X1 U211 ( .IN1(n2508), .IN2(n2570), .IN3(\regf[4][15] ), .IN4(n44), .Q(
        n190) );
  AO22X1 U212 ( .IN1(n2508), .IN2(n2573), .IN3(\regf[4][16] ), .IN4(n44), .Q(
        n191) );
  AO22X1 U213 ( .IN1(n2508), .IN2(n2576), .IN3(\regf[4][17] ), .IN4(n44), .Q(
        n192) );
  AO22X1 U214 ( .IN1(n2509), .IN2(n2579), .IN3(\regf[4][18] ), .IN4(n44), .Q(
        n193) );
  AO22X1 U215 ( .IN1(n2508), .IN2(n2582), .IN3(\regf[4][19] ), .IN4(n44), .Q(
        n194) );
  AO22X1 U216 ( .IN1(n2509), .IN2(n2585), .IN3(\regf[4][20] ), .IN4(n2506), 
        .Q(n195) );
  AO22X1 U217 ( .IN1(n2508), .IN2(n2588), .IN3(\regf[4][21] ), .IN4(n2506), 
        .Q(n196) );
  AO22X1 U218 ( .IN1(n2509), .IN2(n2591), .IN3(\regf[4][22] ), .IN4(n2506), 
        .Q(n197) );
  AO22X1 U219 ( .IN1(n2508), .IN2(n2594), .IN3(\regf[4][23] ), .IN4(n2506), 
        .Q(n198) );
  AO22X1 U220 ( .IN1(n2509), .IN2(n2597), .IN3(\regf[4][24] ), .IN4(n2506), 
        .Q(n199) );
  AO22X1 U221 ( .IN1(n2509), .IN2(n2600), .IN3(\regf[4][25] ), .IN4(n2506), 
        .Q(n200) );
  AO22X1 U222 ( .IN1(n2509), .IN2(n2603), .IN3(\regf[4][26] ), .IN4(n2506), 
        .Q(n201) );
  AO22X1 U223 ( .IN1(n2509), .IN2(n2606), .IN3(\regf[4][27] ), .IN4(n2506), 
        .Q(n202) );
  AO22X1 U224 ( .IN1(n2509), .IN2(n2609), .IN3(\regf[4][28] ), .IN4(n2506), 
        .Q(n203) );
  AO22X1 U225 ( .IN1(n2509), .IN2(n2612), .IN3(\regf[4][29] ), .IN4(n2506), 
        .Q(n204) );
  AO22X1 U226 ( .IN1(n2509), .IN2(n2615), .IN3(\regf[4][30] ), .IN4(n2506), 
        .Q(n205) );
  AO22X1 U227 ( .IN1(n2509), .IN2(n2618), .IN3(\regf[4][31] ), .IN4(n2506), 
        .Q(n206) );
  AO22X1 U228 ( .IN1(n2505), .IN2(n2525), .IN3(\regf[5][0] ), .IN4(n2503), .Q(
        n207) );
  AO22X1 U229 ( .IN1(n2504), .IN2(n2528), .IN3(\regf[5][1] ), .IN4(n2503), .Q(
        n208) );
  AO22X1 U230 ( .IN1(n2505), .IN2(n2531), .IN3(\regf[5][2] ), .IN4(n2503), .Q(
        n209) );
  AO22X1 U231 ( .IN1(n2504), .IN2(n2534), .IN3(\regf[5][3] ), .IN4(n2503), .Q(
        n210) );
  AO22X1 U232 ( .IN1(n2504), .IN2(n2537), .IN3(\regf[5][4] ), .IN4(n2503), .Q(
        n211) );
  AO22X1 U233 ( .IN1(n2505), .IN2(n2540), .IN3(\regf[5][5] ), .IN4(n2503), .Q(
        n212) );
  AO22X1 U234 ( .IN1(n2504), .IN2(n2543), .IN3(\regf[5][6] ), .IN4(n2503), .Q(
        n213) );
  AO22X1 U235 ( .IN1(n2504), .IN2(n2546), .IN3(\regf[5][7] ), .IN4(n2503), .Q(
        n214) );
  AO22X1 U236 ( .IN1(n2505), .IN2(n2549), .IN3(\regf[5][8] ), .IN4(n2503), .Q(
        n215) );
  AO22X1 U237 ( .IN1(n2505), .IN2(n2552), .IN3(\regf[5][9] ), .IN4(n2503), .Q(
        n216) );
  AO22X1 U238 ( .IN1(n2504), .IN2(n2555), .IN3(\regf[5][10] ), .IN4(n2503), 
        .Q(n217) );
  AO22X1 U239 ( .IN1(n2504), .IN2(n2558), .IN3(\regf[5][11] ), .IN4(n2503), 
        .Q(n218) );
  AO22X1 U240 ( .IN1(n2504), .IN2(n2561), .IN3(\regf[5][12] ), .IN4(n2503), 
        .Q(n219) );
  AO22X1 U241 ( .IN1(n2504), .IN2(n2564), .IN3(\regf[5][13] ), .IN4(n2502), 
        .Q(n220) );
  AO22X1 U242 ( .IN1(n2504), .IN2(n2567), .IN3(\regf[5][14] ), .IN4(n46), .Q(
        n221) );
  AO22X1 U243 ( .IN1(n2504), .IN2(n2570), .IN3(\regf[5][15] ), .IN4(n46), .Q(
        n222) );
  AO22X1 U244 ( .IN1(n2504), .IN2(n2573), .IN3(\regf[5][16] ), .IN4(n46), .Q(
        n223) );
  AO22X1 U245 ( .IN1(n2504), .IN2(n2576), .IN3(\regf[5][17] ), .IN4(n46), .Q(
        n224) );
  AO22X1 U246 ( .IN1(n2505), .IN2(n2579), .IN3(\regf[5][18] ), .IN4(n46), .Q(
        n225) );
  AO22X1 U247 ( .IN1(n2504), .IN2(n2582), .IN3(\regf[5][19] ), .IN4(n46), .Q(
        n226) );
  AO22X1 U248 ( .IN1(n2505), .IN2(n2585), .IN3(\regf[5][20] ), .IN4(n2502), 
        .Q(n227) );
  AO22X1 U249 ( .IN1(n2504), .IN2(n2588), .IN3(\regf[5][21] ), .IN4(n2502), 
        .Q(n228) );
  AO22X1 U250 ( .IN1(n2505), .IN2(n2591), .IN3(\regf[5][22] ), .IN4(n2502), 
        .Q(n229) );
  AO22X1 U251 ( .IN1(n2504), .IN2(n2594), .IN3(\regf[5][23] ), .IN4(n2502), 
        .Q(n230) );
  AO22X1 U252 ( .IN1(n2505), .IN2(n2597), .IN3(\regf[5][24] ), .IN4(n2502), 
        .Q(n231) );
  AO22X1 U253 ( .IN1(n2505), .IN2(n2600), .IN3(\regf[5][25] ), .IN4(n2502), 
        .Q(n232) );
  AO22X1 U254 ( .IN1(n2505), .IN2(n2603), .IN3(\regf[5][26] ), .IN4(n2502), 
        .Q(n233) );
  AO22X1 U255 ( .IN1(n2505), .IN2(n2606), .IN3(\regf[5][27] ), .IN4(n2502), 
        .Q(n234) );
  AO22X1 U256 ( .IN1(n2505), .IN2(n2609), .IN3(\regf[5][28] ), .IN4(n2502), 
        .Q(n235) );
  AO22X1 U257 ( .IN1(n2505), .IN2(n2612), .IN3(\regf[5][29] ), .IN4(n2502), 
        .Q(n236) );
  AO22X1 U258 ( .IN1(n2505), .IN2(n2615), .IN3(\regf[5][30] ), .IN4(n2502), 
        .Q(n237) );
  AO22X1 U259 ( .IN1(n2505), .IN2(n2618), .IN3(\regf[5][31] ), .IN4(n2502), 
        .Q(n238) );
  AO22X1 U260 ( .IN1(n2501), .IN2(n2525), .IN3(\regf[6][0] ), .IN4(n2499), .Q(
        n239) );
  AO22X1 U261 ( .IN1(n2500), .IN2(n2528), .IN3(\regf[6][1] ), .IN4(n2499), .Q(
        n240) );
  AO22X1 U262 ( .IN1(n2501), .IN2(n2531), .IN3(\regf[6][2] ), .IN4(n2499), .Q(
        n241) );
  AO22X1 U263 ( .IN1(n2500), .IN2(n2534), .IN3(\regf[6][3] ), .IN4(n2499), .Q(
        n242) );
  AO22X1 U264 ( .IN1(n2500), .IN2(n2537), .IN3(\regf[6][4] ), .IN4(n2499), .Q(
        n243) );
  AO22X1 U265 ( .IN1(n2501), .IN2(n2540), .IN3(\regf[6][5] ), .IN4(n2499), .Q(
        n244) );
  AO22X1 U266 ( .IN1(n2500), .IN2(n2543), .IN3(\regf[6][6] ), .IN4(n2499), .Q(
        n245) );
  AO22X1 U267 ( .IN1(n2500), .IN2(n2546), .IN3(\regf[6][7] ), .IN4(n2499), .Q(
        n246) );
  AO22X1 U268 ( .IN1(n2501), .IN2(n2549), .IN3(\regf[6][8] ), .IN4(n2499), .Q(
        n247) );
  AO22X1 U269 ( .IN1(n2501), .IN2(n2552), .IN3(\regf[6][9] ), .IN4(n2499), .Q(
        n248) );
  AO22X1 U270 ( .IN1(n2500), .IN2(n2555), .IN3(\regf[6][10] ), .IN4(n2499), 
        .Q(n249) );
  AO22X1 U271 ( .IN1(n2500), .IN2(n2558), .IN3(\regf[6][11] ), .IN4(n2499), 
        .Q(n250) );
  AO22X1 U272 ( .IN1(n2500), .IN2(n2561), .IN3(\regf[6][12] ), .IN4(n2499), 
        .Q(n251) );
  AO22X1 U273 ( .IN1(n2500), .IN2(n2564), .IN3(\regf[6][13] ), .IN4(n2498), 
        .Q(n252) );
  AO22X1 U274 ( .IN1(n2500), .IN2(n2567), .IN3(\regf[6][14] ), .IN4(n48), .Q(
        n253) );
  AO22X1 U275 ( .IN1(n2500), .IN2(n2570), .IN3(\regf[6][15] ), .IN4(n48), .Q(
        n254) );
  AO22X1 U276 ( .IN1(n2500), .IN2(n2573), .IN3(\regf[6][16] ), .IN4(n48), .Q(
        n255) );
  AO22X1 U277 ( .IN1(n2500), .IN2(n2576), .IN3(\regf[6][17] ), .IN4(n48), .Q(
        n256) );
  AO22X1 U278 ( .IN1(n2501), .IN2(n2579), .IN3(\regf[6][18] ), .IN4(n48), .Q(
        n257) );
  AO22X1 U279 ( .IN1(n2500), .IN2(n2582), .IN3(\regf[6][19] ), .IN4(n48), .Q(
        n258) );
  AO22X1 U280 ( .IN1(n2501), .IN2(n2585), .IN3(\regf[6][20] ), .IN4(n2498), 
        .Q(n259) );
  AO22X1 U281 ( .IN1(n2500), .IN2(n2588), .IN3(\regf[6][21] ), .IN4(n2498), 
        .Q(n260) );
  AO22X1 U282 ( .IN1(n2501), .IN2(n2591), .IN3(\regf[6][22] ), .IN4(n2498), 
        .Q(n261) );
  AO22X1 U283 ( .IN1(n2500), .IN2(n2594), .IN3(\regf[6][23] ), .IN4(n2498), 
        .Q(n262) );
  AO22X1 U284 ( .IN1(n2501), .IN2(n2597), .IN3(\regf[6][24] ), .IN4(n2498), 
        .Q(n263) );
  AO22X1 U285 ( .IN1(n2501), .IN2(n2600), .IN3(\regf[6][25] ), .IN4(n2498), 
        .Q(n264) );
  AO22X1 U286 ( .IN1(n2501), .IN2(n2603), .IN3(\regf[6][26] ), .IN4(n2498), 
        .Q(n265) );
  AO22X1 U287 ( .IN1(n2501), .IN2(n2606), .IN3(\regf[6][27] ), .IN4(n2498), 
        .Q(n266) );
  AO22X1 U288 ( .IN1(n2501), .IN2(n2609), .IN3(\regf[6][28] ), .IN4(n2498), 
        .Q(n267) );
  AO22X1 U289 ( .IN1(n2501), .IN2(n2612), .IN3(\regf[6][29] ), .IN4(n2498), 
        .Q(n268) );
  AO22X1 U290 ( .IN1(n2501), .IN2(n2615), .IN3(\regf[6][30] ), .IN4(n2498), 
        .Q(n269) );
  AO22X1 U291 ( .IN1(n2501), .IN2(n2618), .IN3(\regf[6][31] ), .IN4(n2498), 
        .Q(n270) );
  AO22X1 U292 ( .IN1(n2497), .IN2(n2525), .IN3(\regf[7][0] ), .IN4(n2495), .Q(
        n271) );
  AO22X1 U293 ( .IN1(n2496), .IN2(n2528), .IN3(\regf[7][1] ), .IN4(n2495), .Q(
        n272) );
  AO22X1 U294 ( .IN1(n2497), .IN2(n2531), .IN3(\regf[7][2] ), .IN4(n2495), .Q(
        n273) );
  AO22X1 U295 ( .IN1(n2496), .IN2(n2534), .IN3(\regf[7][3] ), .IN4(n2495), .Q(
        n274) );
  AO22X1 U296 ( .IN1(n2496), .IN2(n2537), .IN3(\regf[7][4] ), .IN4(n2495), .Q(
        n275) );
  AO22X1 U297 ( .IN1(n2497), .IN2(n2540), .IN3(\regf[7][5] ), .IN4(n2495), .Q(
        n276) );
  AO22X1 U298 ( .IN1(n2496), .IN2(n2543), .IN3(\regf[7][6] ), .IN4(n2495), .Q(
        n277) );
  AO22X1 U299 ( .IN1(n2496), .IN2(n2546), .IN3(\regf[7][7] ), .IN4(n2495), .Q(
        n278) );
  AO22X1 U300 ( .IN1(n2497), .IN2(n2549), .IN3(\regf[7][8] ), .IN4(n2495), .Q(
        n279) );
  AO22X1 U301 ( .IN1(n2497), .IN2(n2552), .IN3(\regf[7][9] ), .IN4(n2495), .Q(
        n280) );
  AO22X1 U302 ( .IN1(n2496), .IN2(n2555), .IN3(\regf[7][10] ), .IN4(n2495), 
        .Q(n281) );
  AO22X1 U303 ( .IN1(n2496), .IN2(n2558), .IN3(\regf[7][11] ), .IN4(n2495), 
        .Q(n282) );
  AO22X1 U304 ( .IN1(n2496), .IN2(n2561), .IN3(\regf[7][12] ), .IN4(n2495), 
        .Q(n283) );
  AO22X1 U305 ( .IN1(n2496), .IN2(n2564), .IN3(\regf[7][13] ), .IN4(n2494), 
        .Q(n284) );
  AO22X1 U306 ( .IN1(n2496), .IN2(n2567), .IN3(\regf[7][14] ), .IN4(n50), .Q(
        n285) );
  AO22X1 U307 ( .IN1(n2496), .IN2(n2570), .IN3(\regf[7][15] ), .IN4(n50), .Q(
        n286) );
  AO22X1 U308 ( .IN1(n2496), .IN2(n2573), .IN3(\regf[7][16] ), .IN4(n50), .Q(
        n287) );
  AO22X1 U309 ( .IN1(n2496), .IN2(n2576), .IN3(\regf[7][17] ), .IN4(n50), .Q(
        n288) );
  AO22X1 U310 ( .IN1(n2497), .IN2(n2579), .IN3(\regf[7][18] ), .IN4(n50), .Q(
        n289) );
  AO22X1 U311 ( .IN1(n2496), .IN2(n2582), .IN3(\regf[7][19] ), .IN4(n50), .Q(
        n290) );
  AO22X1 U312 ( .IN1(n2497), .IN2(n2585), .IN3(\regf[7][20] ), .IN4(n2494), 
        .Q(n291) );
  AO22X1 U313 ( .IN1(n2496), .IN2(n2588), .IN3(\regf[7][21] ), .IN4(n2494), 
        .Q(n292) );
  AO22X1 U314 ( .IN1(n2497), .IN2(n2591), .IN3(\regf[7][22] ), .IN4(n2494), 
        .Q(n293) );
  AO22X1 U315 ( .IN1(n2496), .IN2(n2594), .IN3(\regf[7][23] ), .IN4(n2494), 
        .Q(n294) );
  AO22X1 U316 ( .IN1(n2497), .IN2(n2597), .IN3(\regf[7][24] ), .IN4(n2494), 
        .Q(n295) );
  AO22X1 U317 ( .IN1(n2497), .IN2(n2600), .IN3(\regf[7][25] ), .IN4(n2494), 
        .Q(n296) );
  AO22X1 U318 ( .IN1(n2497), .IN2(n2603), .IN3(\regf[7][26] ), .IN4(n2494), 
        .Q(n297) );
  AO22X1 U319 ( .IN1(n2497), .IN2(n2606), .IN3(\regf[7][27] ), .IN4(n2494), 
        .Q(n298) );
  AO22X1 U320 ( .IN1(n2497), .IN2(n2609), .IN3(\regf[7][28] ), .IN4(n2494), 
        .Q(n299) );
  AO22X1 U321 ( .IN1(n2497), .IN2(n2612), .IN3(\regf[7][29] ), .IN4(n2494), 
        .Q(n300) );
  AO22X1 U322 ( .IN1(n2497), .IN2(n2615), .IN3(\regf[7][30] ), .IN4(n2494), 
        .Q(n301) );
  AO22X1 U323 ( .IN1(n2497), .IN2(n2618), .IN3(\regf[7][31] ), .IN4(n2494), 
        .Q(n302) );
  AND3X1 U324 ( .IN1(n2712), .IN2(n2711), .IN3(wr_en), .Q(n39) );
  AO22X1 U325 ( .IN1(n2493), .IN2(n2525), .IN3(\regf[8][0] ), .IN4(n2491), .Q(
        n303) );
  AO22X1 U326 ( .IN1(n2492), .IN2(n2528), .IN3(\regf[8][1] ), .IN4(n2491), .Q(
        n304) );
  AO22X1 U327 ( .IN1(n2493), .IN2(n2531), .IN3(\regf[8][2] ), .IN4(n2491), .Q(
        n305) );
  AO22X1 U328 ( .IN1(n2492), .IN2(n2534), .IN3(\regf[8][3] ), .IN4(n2491), .Q(
        n306) );
  AO22X1 U329 ( .IN1(n2493), .IN2(n2537), .IN3(\regf[8][4] ), .IN4(n2491), .Q(
        n307) );
  AO22X1 U330 ( .IN1(n2492), .IN2(n2540), .IN3(\regf[8][5] ), .IN4(n2491), .Q(
        n308) );
  AO22X1 U331 ( .IN1(n2492), .IN2(n2543), .IN3(\regf[8][6] ), .IN4(n2491), .Q(
        n309) );
  AO22X1 U332 ( .IN1(n2493), .IN2(n2546), .IN3(\regf[8][7] ), .IN4(n2491), .Q(
        n310) );
  AO22X1 U333 ( .IN1(n2492), .IN2(n2549), .IN3(\regf[8][8] ), .IN4(n2491), .Q(
        n311) );
  AO22X1 U334 ( .IN1(n2492), .IN2(n2552), .IN3(\regf[8][9] ), .IN4(n2491), .Q(
        n312) );
  AO22X1 U335 ( .IN1(n2493), .IN2(n2555), .IN3(\regf[8][10] ), .IN4(n2491), 
        .Q(n313) );
  AO22X1 U336 ( .IN1(n2493), .IN2(n2558), .IN3(\regf[8][11] ), .IN4(n2491), 
        .Q(n314) );
  AO22X1 U337 ( .IN1(n2492), .IN2(n2561), .IN3(\regf[8][12] ), .IN4(n2491), 
        .Q(n315) );
  AO22X1 U338 ( .IN1(n2493), .IN2(n2564), .IN3(\regf[8][13] ), .IN4(n2490), 
        .Q(n316) );
  AO22X1 U339 ( .IN1(n2492), .IN2(n2567), .IN3(\regf[8][14] ), .IN4(n52), .Q(
        n317) );
  AO22X1 U340 ( .IN1(n2493), .IN2(n2570), .IN3(\regf[8][15] ), .IN4(n52), .Q(
        n318) );
  AO22X1 U341 ( .IN1(n2492), .IN2(n2573), .IN3(\regf[8][16] ), .IN4(n52), .Q(
        n319) );
  AO22X1 U342 ( .IN1(n2493), .IN2(n2576), .IN3(\regf[8][17] ), .IN4(n52), .Q(
        n320) );
  AO22X1 U343 ( .IN1(n2492), .IN2(n2579), .IN3(\regf[8][18] ), .IN4(n52), .Q(
        n321) );
  AO22X1 U344 ( .IN1(n2492), .IN2(n2582), .IN3(\regf[8][19] ), .IN4(n52), .Q(
        n322) );
  AO22X1 U345 ( .IN1(n2492), .IN2(n2585), .IN3(\regf[8][20] ), .IN4(n2490), 
        .Q(n323) );
  AO22X1 U346 ( .IN1(n2492), .IN2(n2588), .IN3(\regf[8][21] ), .IN4(n2490), 
        .Q(n324) );
  AO22X1 U347 ( .IN1(n2492), .IN2(n2591), .IN3(\regf[8][22] ), .IN4(n2490), 
        .Q(n325) );
  AO22X1 U348 ( .IN1(n2492), .IN2(n2594), .IN3(\regf[8][23] ), .IN4(n2490), 
        .Q(n326) );
  AO22X1 U349 ( .IN1(n2492), .IN2(n2597), .IN3(\regf[8][24] ), .IN4(n2490), 
        .Q(n327) );
  AO22X1 U350 ( .IN1(n2493), .IN2(n2600), .IN3(\regf[8][25] ), .IN4(n2490), 
        .Q(n328) );
  AO22X1 U351 ( .IN1(n2493), .IN2(n2603), .IN3(\regf[8][26] ), .IN4(n2490), 
        .Q(n329) );
  AO22X1 U352 ( .IN1(n2493), .IN2(n2606), .IN3(\regf[8][27] ), .IN4(n2490), 
        .Q(n330) );
  AO22X1 U353 ( .IN1(n2493), .IN2(n2609), .IN3(\regf[8][28] ), .IN4(n2490), 
        .Q(n331) );
  AO22X1 U354 ( .IN1(n2493), .IN2(n2612), .IN3(\regf[8][29] ), .IN4(n2490), 
        .Q(n332) );
  AO22X1 U355 ( .IN1(n2493), .IN2(n2615), .IN3(\regf[8][30] ), .IN4(n2490), 
        .Q(n333) );
  AO22X1 U356 ( .IN1(n2493), .IN2(n2618), .IN3(\regf[8][31] ), .IN4(n2490), 
        .Q(n334) );
  AO22X1 U357 ( .IN1(n2487), .IN2(n2525), .IN3(\regf[9][0] ), .IN4(n2486), .Q(
        n335) );
  AO22X1 U358 ( .IN1(n2487), .IN2(n2528), .IN3(\regf[9][1] ), .IN4(n2486), .Q(
        n336) );
  AO22X1 U359 ( .IN1(n2487), .IN2(n2531), .IN3(\regf[9][2] ), .IN4(n2486), .Q(
        n337) );
  AO22X1 U360 ( .IN1(n2487), .IN2(n2534), .IN3(\regf[9][3] ), .IN4(n2486), .Q(
        n338) );
  AO22X1 U361 ( .IN1(n2488), .IN2(n2537), .IN3(\regf[9][4] ), .IN4(n2486), .Q(
        n339) );
  AO22X1 U362 ( .IN1(n2489), .IN2(n2540), .IN3(\regf[9][5] ), .IN4(n2486), .Q(
        n340) );
  AO22X1 U363 ( .IN1(n2488), .IN2(n2543), .IN3(\regf[9][6] ), .IN4(n2486), .Q(
        n341) );
  AO22X1 U364 ( .IN1(n2488), .IN2(n2546), .IN3(\regf[9][7] ), .IN4(n2486), .Q(
        n342) );
  AO22X1 U365 ( .IN1(n2489), .IN2(n2549), .IN3(\regf[9][8] ), .IN4(n2486), .Q(
        n343) );
  AO22X1 U366 ( .IN1(n2489), .IN2(n2552), .IN3(\regf[9][9] ), .IN4(n2486), .Q(
        n344) );
  AO22X1 U367 ( .IN1(n2488), .IN2(n2555), .IN3(\regf[9][10] ), .IN4(n2486), 
        .Q(n345) );
  AO22X1 U368 ( .IN1(n2488), .IN2(n2558), .IN3(\regf[9][11] ), .IN4(n2486), 
        .Q(n346) );
  AO22X1 U369 ( .IN1(n2488), .IN2(n2561), .IN3(\regf[9][12] ), .IN4(n2486), 
        .Q(n347) );
  AO22X1 U370 ( .IN1(n2488), .IN2(n2564), .IN3(\regf[9][13] ), .IN4(n2485), 
        .Q(n348) );
  AO22X1 U371 ( .IN1(n2488), .IN2(n2567), .IN3(\regf[9][14] ), .IN4(n54), .Q(
        n349) );
  AO22X1 U372 ( .IN1(n2488), .IN2(n2570), .IN3(\regf[9][15] ), .IN4(n54), .Q(
        n350) );
  AO22X1 U373 ( .IN1(n2488), .IN2(n2573), .IN3(\regf[9][16] ), .IN4(n54), .Q(
        n351) );
  AO22X1 U374 ( .IN1(n2488), .IN2(n2576), .IN3(\regf[9][17] ), .IN4(n54), .Q(
        n352) );
  AO22X1 U375 ( .IN1(n2489), .IN2(n2579), .IN3(\regf[9][18] ), .IN4(n54), .Q(
        n353) );
  AO22X1 U376 ( .IN1(n2488), .IN2(n2582), .IN3(\regf[9][19] ), .IN4(n54), .Q(
        n354) );
  AO22X1 U377 ( .IN1(n2489), .IN2(n2585), .IN3(\regf[9][20] ), .IN4(n2485), 
        .Q(n355) );
  AO22X1 U378 ( .IN1(n2488), .IN2(n2588), .IN3(\regf[9][21] ), .IN4(n2485), 
        .Q(n356) );
  AO22X1 U379 ( .IN1(n2489), .IN2(n2591), .IN3(\regf[9][22] ), .IN4(n2485), 
        .Q(n357) );
  AO22X1 U380 ( .IN1(n2488), .IN2(n2594), .IN3(\regf[9][23] ), .IN4(n2485), 
        .Q(n358) );
  AO22X1 U381 ( .IN1(n2489), .IN2(n2597), .IN3(\regf[9][24] ), .IN4(n2485), 
        .Q(n359) );
  AO22X1 U382 ( .IN1(n2489), .IN2(n2600), .IN3(\regf[9][25] ), .IN4(n2485), 
        .Q(n360) );
  AO22X1 U383 ( .IN1(n2489), .IN2(n2603), .IN3(\regf[9][26] ), .IN4(n2485), 
        .Q(n361) );
  AO22X1 U384 ( .IN1(n2489), .IN2(n2606), .IN3(\regf[9][27] ), .IN4(n2485), 
        .Q(n362) );
  AO22X1 U385 ( .IN1(n2489), .IN2(n2609), .IN3(\regf[9][28] ), .IN4(n2485), 
        .Q(n363) );
  AO22X1 U386 ( .IN1(n2489), .IN2(n2612), .IN3(\regf[9][29] ), .IN4(n2485), 
        .Q(n364) );
  AO22X1 U387 ( .IN1(n2489), .IN2(n2615), .IN3(\regf[9][30] ), .IN4(n2485), 
        .Q(n365) );
  AO22X1 U388 ( .IN1(n2489), .IN2(n2618), .IN3(\regf[9][31] ), .IN4(n2485), 
        .Q(n366) );
  AO22X1 U389 ( .IN1(n2482), .IN2(n2525), .IN3(\regf[10][0] ), .IN4(n2481), 
        .Q(n367) );
  AO22X1 U390 ( .IN1(n2482), .IN2(n2528), .IN3(\regf[10][1] ), .IN4(n2481), 
        .Q(n368) );
  AO22X1 U391 ( .IN1(n2482), .IN2(n2531), .IN3(\regf[10][2] ), .IN4(n2481), 
        .Q(n369) );
  AO22X1 U392 ( .IN1(n2482), .IN2(n2534), .IN3(\regf[10][3] ), .IN4(n2481), 
        .Q(n370) );
  AO22X1 U393 ( .IN1(n2483), .IN2(n2537), .IN3(\regf[10][4] ), .IN4(n2481), 
        .Q(n371) );
  AO22X1 U394 ( .IN1(n2484), .IN2(n2540), .IN3(\regf[10][5] ), .IN4(n2481), 
        .Q(n372) );
  AO22X1 U395 ( .IN1(n2483), .IN2(n2543), .IN3(\regf[10][6] ), .IN4(n2481), 
        .Q(n373) );
  AO22X1 U396 ( .IN1(n2483), .IN2(n2546), .IN3(\regf[10][7] ), .IN4(n2481), 
        .Q(n374) );
  AO22X1 U397 ( .IN1(n2484), .IN2(n2549), .IN3(\regf[10][8] ), .IN4(n2481), 
        .Q(n375) );
  AO22X1 U398 ( .IN1(n2484), .IN2(n2552), .IN3(\regf[10][9] ), .IN4(n2481), 
        .Q(n376) );
  AO22X1 U399 ( .IN1(n2483), .IN2(n2555), .IN3(\regf[10][10] ), .IN4(n2481), 
        .Q(n377) );
  AO22X1 U400 ( .IN1(n2483), .IN2(n2558), .IN3(\regf[10][11] ), .IN4(n2481), 
        .Q(n378) );
  AO22X1 U401 ( .IN1(n2483), .IN2(n2561), .IN3(\regf[10][12] ), .IN4(n2481), 
        .Q(n379) );
  AO22X1 U402 ( .IN1(n2483), .IN2(n2564), .IN3(\regf[10][13] ), .IN4(n2480), 
        .Q(n380) );
  AO22X1 U403 ( .IN1(n2483), .IN2(n2567), .IN3(\regf[10][14] ), .IN4(n55), .Q(
        n381) );
  AO22X1 U404 ( .IN1(n2483), .IN2(n2570), .IN3(\regf[10][15] ), .IN4(n55), .Q(
        n382) );
  AO22X1 U405 ( .IN1(n2483), .IN2(n2573), .IN3(\regf[10][16] ), .IN4(n55), .Q(
        n383) );
  AO22X1 U406 ( .IN1(n2483), .IN2(n2576), .IN3(\regf[10][17] ), .IN4(n55), .Q(
        n384) );
  AO22X1 U407 ( .IN1(n2484), .IN2(n2579), .IN3(\regf[10][18] ), .IN4(n55), .Q(
        n385) );
  AO22X1 U408 ( .IN1(n2483), .IN2(n2582), .IN3(\regf[10][19] ), .IN4(n55), .Q(
        n386) );
  AO22X1 U409 ( .IN1(n2484), .IN2(n2585), .IN3(\regf[10][20] ), .IN4(n2480), 
        .Q(n387) );
  AO22X1 U410 ( .IN1(n2483), .IN2(n2588), .IN3(\regf[10][21] ), .IN4(n2480), 
        .Q(n388) );
  AO22X1 U411 ( .IN1(n2484), .IN2(n2591), .IN3(\regf[10][22] ), .IN4(n2480), 
        .Q(n389) );
  AO22X1 U412 ( .IN1(n2483), .IN2(n2594), .IN3(\regf[10][23] ), .IN4(n2480), 
        .Q(n390) );
  AO22X1 U413 ( .IN1(n2484), .IN2(n2597), .IN3(\regf[10][24] ), .IN4(n2480), 
        .Q(n391) );
  AO22X1 U414 ( .IN1(n2484), .IN2(n2600), .IN3(\regf[10][25] ), .IN4(n2480), 
        .Q(n392) );
  AO22X1 U415 ( .IN1(n2484), .IN2(n2603), .IN3(\regf[10][26] ), .IN4(n2480), 
        .Q(n393) );
  AO22X1 U416 ( .IN1(n2484), .IN2(n2606), .IN3(\regf[10][27] ), .IN4(n2480), 
        .Q(n394) );
  AO22X1 U417 ( .IN1(n2484), .IN2(n2609), .IN3(\regf[10][28] ), .IN4(n2480), 
        .Q(n395) );
  AO22X1 U418 ( .IN1(n2484), .IN2(n2612), .IN3(\regf[10][29] ), .IN4(n2480), 
        .Q(n396) );
  AO22X1 U419 ( .IN1(n2484), .IN2(n2615), .IN3(\regf[10][30] ), .IN4(n2480), 
        .Q(n397) );
  AO22X1 U420 ( .IN1(n2484), .IN2(n2618), .IN3(\regf[10][31] ), .IN4(n2480), 
        .Q(n398) );
  AO22X1 U421 ( .IN1(n2477), .IN2(n2525), .IN3(\regf[11][0] ), .IN4(n2476), 
        .Q(n399) );
  AO22X1 U422 ( .IN1(n2477), .IN2(n2528), .IN3(\regf[11][1] ), .IN4(n2476), 
        .Q(n400) );
  AO22X1 U423 ( .IN1(n2477), .IN2(n2531), .IN3(\regf[11][2] ), .IN4(n2476), 
        .Q(n401) );
  AO22X1 U424 ( .IN1(n2477), .IN2(n2534), .IN3(\regf[11][3] ), .IN4(n2476), 
        .Q(n402) );
  AO22X1 U425 ( .IN1(n2479), .IN2(n2537), .IN3(\regf[11][4] ), .IN4(n2476), 
        .Q(n403) );
  AO22X1 U426 ( .IN1(n2478), .IN2(n2540), .IN3(\regf[11][5] ), .IN4(n2476), 
        .Q(n404) );
  AO22X1 U427 ( .IN1(n2478), .IN2(n2543), .IN3(\regf[11][6] ), .IN4(n2476), 
        .Q(n405) );
  AO22X1 U428 ( .IN1(n2479), .IN2(n2546), .IN3(\regf[11][7] ), .IN4(n2476), 
        .Q(n406) );
  AO22X1 U429 ( .IN1(n2478), .IN2(n2549), .IN3(\regf[11][8] ), .IN4(n2476), 
        .Q(n407) );
  AO22X1 U430 ( .IN1(n2478), .IN2(n2552), .IN3(\regf[11][9] ), .IN4(n2476), 
        .Q(n408) );
  AO22X1 U431 ( .IN1(n2479), .IN2(n2555), .IN3(\regf[11][10] ), .IN4(n2476), 
        .Q(n409) );
  AO22X1 U432 ( .IN1(n2479), .IN2(n2558), .IN3(\regf[11][11] ), .IN4(n2476), 
        .Q(n410) );
  AO22X1 U433 ( .IN1(n2478), .IN2(n2561), .IN3(\regf[11][12] ), .IN4(n2476), 
        .Q(n411) );
  AO22X1 U434 ( .IN1(n2479), .IN2(n2564), .IN3(\regf[11][13] ), .IN4(n2475), 
        .Q(n412) );
  AO22X1 U435 ( .IN1(n2478), .IN2(n2567), .IN3(\regf[11][14] ), .IN4(n56), .Q(
        n413) );
  AO22X1 U436 ( .IN1(n2479), .IN2(n2570), .IN3(\regf[11][15] ), .IN4(n56), .Q(
        n414) );
  AO22X1 U437 ( .IN1(n2478), .IN2(n2573), .IN3(\regf[11][16] ), .IN4(n56), .Q(
        n415) );
  AO22X1 U438 ( .IN1(n2479), .IN2(n2576), .IN3(\regf[11][17] ), .IN4(n56), .Q(
        n416) );
  AO22X1 U439 ( .IN1(n2478), .IN2(n2579), .IN3(\regf[11][18] ), .IN4(n56), .Q(
        n417) );
  AO22X1 U440 ( .IN1(n2478), .IN2(n2582), .IN3(\regf[11][19] ), .IN4(n56), .Q(
        n418) );
  AO22X1 U441 ( .IN1(n2478), .IN2(n2585), .IN3(\regf[11][20] ), .IN4(n2475), 
        .Q(n419) );
  AO22X1 U442 ( .IN1(n2478), .IN2(n2588), .IN3(\regf[11][21] ), .IN4(n2475), 
        .Q(n420) );
  AO22X1 U443 ( .IN1(n2478), .IN2(n2591), .IN3(\regf[11][22] ), .IN4(n2475), 
        .Q(n421) );
  AO22X1 U444 ( .IN1(n2478), .IN2(n2594), .IN3(\regf[11][23] ), .IN4(n2475), 
        .Q(n422) );
  AO22X1 U445 ( .IN1(n2478), .IN2(n2597), .IN3(\regf[11][24] ), .IN4(n2475), 
        .Q(n423) );
  AO22X1 U446 ( .IN1(n2479), .IN2(n2600), .IN3(\regf[11][25] ), .IN4(n2475), 
        .Q(n424) );
  AO22X1 U447 ( .IN1(n2479), .IN2(n2603), .IN3(\regf[11][26] ), .IN4(n2475), 
        .Q(n425) );
  AO22X1 U448 ( .IN1(n2479), .IN2(n2606), .IN3(\regf[11][27] ), .IN4(n2475), 
        .Q(n426) );
  AO22X1 U449 ( .IN1(n2479), .IN2(n2609), .IN3(\regf[11][28] ), .IN4(n2475), 
        .Q(n427) );
  AO22X1 U450 ( .IN1(n2479), .IN2(n2612), .IN3(\regf[11][29] ), .IN4(n2475), 
        .Q(n428) );
  AO22X1 U451 ( .IN1(n2479), .IN2(n2615), .IN3(\regf[11][30] ), .IN4(n2475), 
        .Q(n429) );
  AO22X1 U452 ( .IN1(n2479), .IN2(n2618), .IN3(\regf[11][31] ), .IN4(n2475), 
        .Q(n430) );
  AO22X1 U453 ( .IN1(n2474), .IN2(n2525), .IN3(\regf[12][0] ), .IN4(n2472), 
        .Q(n431) );
  AO22X1 U454 ( .IN1(n2473), .IN2(n2528), .IN3(\regf[12][1] ), .IN4(n2472), 
        .Q(n432) );
  AO22X1 U455 ( .IN1(n2474), .IN2(n2531), .IN3(\regf[12][2] ), .IN4(n2472), 
        .Q(n433) );
  AO22X1 U456 ( .IN1(n2473), .IN2(n2534), .IN3(\regf[12][3] ), .IN4(n2472), 
        .Q(n434) );
  AO22X1 U457 ( .IN1(n2473), .IN2(n2537), .IN3(\regf[12][4] ), .IN4(n2472), 
        .Q(n435) );
  AO22X1 U458 ( .IN1(n2474), .IN2(n2540), .IN3(\regf[12][5] ), .IN4(n2472), 
        .Q(n436) );
  AO22X1 U459 ( .IN1(n2473), .IN2(n2543), .IN3(\regf[12][6] ), .IN4(n2472), 
        .Q(n437) );
  AO22X1 U460 ( .IN1(n2473), .IN2(n2546), .IN3(\regf[12][7] ), .IN4(n2472), 
        .Q(n438) );
  AO22X1 U461 ( .IN1(n2474), .IN2(n2549), .IN3(\regf[12][8] ), .IN4(n2472), 
        .Q(n439) );
  AO22X1 U462 ( .IN1(n2474), .IN2(n2552), .IN3(\regf[12][9] ), .IN4(n2472), 
        .Q(n440) );
  AO22X1 U463 ( .IN1(n2473), .IN2(n2555), .IN3(\regf[12][10] ), .IN4(n2472), 
        .Q(n441) );
  AO22X1 U464 ( .IN1(n2473), .IN2(n2558), .IN3(\regf[12][11] ), .IN4(n2472), 
        .Q(n442) );
  AO22X1 U465 ( .IN1(n2473), .IN2(n2561), .IN3(\regf[12][12] ), .IN4(n2472), 
        .Q(n443) );
  AO22X1 U466 ( .IN1(n2473), .IN2(n2564), .IN3(\regf[12][13] ), .IN4(n2471), 
        .Q(n444) );
  AO22X1 U467 ( .IN1(n2473), .IN2(n2567), .IN3(\regf[12][14] ), .IN4(n57), .Q(
        n445) );
  AO22X1 U468 ( .IN1(n2473), .IN2(n2570), .IN3(\regf[12][15] ), .IN4(n57), .Q(
        n446) );
  AO22X1 U469 ( .IN1(n2473), .IN2(n2573), .IN3(\regf[12][16] ), .IN4(n57), .Q(
        n447) );
  AO22X1 U470 ( .IN1(n2473), .IN2(n2576), .IN3(\regf[12][17] ), .IN4(n57), .Q(
        n448) );
  AO22X1 U471 ( .IN1(n2474), .IN2(n2579), .IN3(\regf[12][18] ), .IN4(n57), .Q(
        n449) );
  AO22X1 U472 ( .IN1(n2473), .IN2(n2582), .IN3(\regf[12][19] ), .IN4(n57), .Q(
        n450) );
  AO22X1 U473 ( .IN1(n2474), .IN2(n2585), .IN3(\regf[12][20] ), .IN4(n2471), 
        .Q(n451) );
  AO22X1 U474 ( .IN1(n2473), .IN2(n2588), .IN3(\regf[12][21] ), .IN4(n2471), 
        .Q(n452) );
  AO22X1 U475 ( .IN1(n2474), .IN2(n2591), .IN3(\regf[12][22] ), .IN4(n2471), 
        .Q(n453) );
  AO22X1 U476 ( .IN1(n2473), .IN2(n2594), .IN3(\regf[12][23] ), .IN4(n2471), 
        .Q(n454) );
  AO22X1 U477 ( .IN1(n2474), .IN2(n2597), .IN3(\regf[12][24] ), .IN4(n2471), 
        .Q(n455) );
  AO22X1 U478 ( .IN1(n2474), .IN2(n2600), .IN3(\regf[12][25] ), .IN4(n2471), 
        .Q(n456) );
  AO22X1 U479 ( .IN1(n2474), .IN2(n2603), .IN3(\regf[12][26] ), .IN4(n2471), 
        .Q(n457) );
  AO22X1 U480 ( .IN1(n2474), .IN2(n2606), .IN3(\regf[12][27] ), .IN4(n2471), 
        .Q(n458) );
  AO22X1 U481 ( .IN1(n2474), .IN2(n2609), .IN3(\regf[12][28] ), .IN4(n2471), 
        .Q(n459) );
  AO22X1 U482 ( .IN1(n2474), .IN2(n2612), .IN3(\regf[12][29] ), .IN4(n2471), 
        .Q(n460) );
  AO22X1 U483 ( .IN1(n2474), .IN2(n2615), .IN3(\regf[12][30] ), .IN4(n2471), 
        .Q(n461) );
  AO22X1 U484 ( .IN1(n2474), .IN2(n2618), .IN3(\regf[12][31] ), .IN4(n2471), 
        .Q(n462) );
  AO22X1 U485 ( .IN1(n2470), .IN2(n2526), .IN3(\regf[13][0] ), .IN4(n2468), 
        .Q(n463) );
  AO22X1 U486 ( .IN1(n2469), .IN2(n2529), .IN3(\regf[13][1] ), .IN4(n2468), 
        .Q(n464) );
  AO22X1 U487 ( .IN1(n2470), .IN2(n2532), .IN3(\regf[13][2] ), .IN4(n2468), 
        .Q(n465) );
  AO22X1 U488 ( .IN1(n2469), .IN2(n2535), .IN3(\regf[13][3] ), .IN4(n2468), 
        .Q(n466) );
  AO22X1 U489 ( .IN1(n2469), .IN2(n2538), .IN3(\regf[13][4] ), .IN4(n2468), 
        .Q(n467) );
  AO22X1 U490 ( .IN1(n2470), .IN2(n2541), .IN3(\regf[13][5] ), .IN4(n2468), 
        .Q(n468) );
  AO22X1 U491 ( .IN1(n2469), .IN2(n2544), .IN3(\regf[13][6] ), .IN4(n2468), 
        .Q(n469) );
  AO22X1 U492 ( .IN1(n2469), .IN2(n2547), .IN3(\regf[13][7] ), .IN4(n2468), 
        .Q(n470) );
  AO22X1 U493 ( .IN1(n2470), .IN2(n2550), .IN3(\regf[13][8] ), .IN4(n2468), 
        .Q(n471) );
  AO22X1 U494 ( .IN1(n2470), .IN2(n2553), .IN3(\regf[13][9] ), .IN4(n2468), 
        .Q(n472) );
  AO22X1 U495 ( .IN1(n2469), .IN2(n2556), .IN3(\regf[13][10] ), .IN4(n2468), 
        .Q(n473) );
  AO22X1 U496 ( .IN1(n2469), .IN2(n2559), .IN3(\regf[13][11] ), .IN4(n2468), 
        .Q(n474) );
  AO22X1 U497 ( .IN1(n2469), .IN2(n2562), .IN3(\regf[13][12] ), .IN4(n2468), 
        .Q(n475) );
  AO22X1 U498 ( .IN1(n2469), .IN2(n2565), .IN3(\regf[13][13] ), .IN4(n2467), 
        .Q(n476) );
  AO22X1 U499 ( .IN1(n2469), .IN2(n2568), .IN3(\regf[13][14] ), .IN4(n58), .Q(
        n477) );
  AO22X1 U500 ( .IN1(n2469), .IN2(n2571), .IN3(\regf[13][15] ), .IN4(n58), .Q(
        n478) );
  AO22X1 U501 ( .IN1(n2469), .IN2(n2574), .IN3(\regf[13][16] ), .IN4(n58), .Q(
        n479) );
  AO22X1 U502 ( .IN1(n2469), .IN2(n2577), .IN3(\regf[13][17] ), .IN4(n58), .Q(
        n480) );
  AO22X1 U503 ( .IN1(n2470), .IN2(n2580), .IN3(\regf[13][18] ), .IN4(n58), .Q(
        n481) );
  AO22X1 U504 ( .IN1(n2469), .IN2(n2583), .IN3(\regf[13][19] ), .IN4(n58), .Q(
        n482) );
  AO22X1 U505 ( .IN1(n2470), .IN2(n2586), .IN3(\regf[13][20] ), .IN4(n2467), 
        .Q(n483) );
  AO22X1 U506 ( .IN1(n2469), .IN2(n2589), .IN3(\regf[13][21] ), .IN4(n2467), 
        .Q(n484) );
  AO22X1 U507 ( .IN1(n2470), .IN2(n2592), .IN3(\regf[13][22] ), .IN4(n2467), 
        .Q(n485) );
  AO22X1 U508 ( .IN1(n2469), .IN2(n2595), .IN3(\regf[13][23] ), .IN4(n2467), 
        .Q(n486) );
  AO22X1 U509 ( .IN1(n2470), .IN2(n2598), .IN3(\regf[13][24] ), .IN4(n2467), 
        .Q(n487) );
  AO22X1 U510 ( .IN1(n2470), .IN2(n2601), .IN3(\regf[13][25] ), .IN4(n2467), 
        .Q(n488) );
  AO22X1 U511 ( .IN1(n2470), .IN2(n2604), .IN3(\regf[13][26] ), .IN4(n2467), 
        .Q(n489) );
  AO22X1 U512 ( .IN1(n2470), .IN2(n2607), .IN3(\regf[13][27] ), .IN4(n2467), 
        .Q(n490) );
  AO22X1 U513 ( .IN1(n2470), .IN2(n2610), .IN3(\regf[13][28] ), .IN4(n2467), 
        .Q(n491) );
  AO22X1 U514 ( .IN1(n2470), .IN2(n2613), .IN3(\regf[13][29] ), .IN4(n2467), 
        .Q(n492) );
  AO22X1 U515 ( .IN1(n2470), .IN2(n2616), .IN3(\regf[13][30] ), .IN4(n2467), 
        .Q(n493) );
  AO22X1 U516 ( .IN1(n2470), .IN2(n2619), .IN3(\regf[13][31] ), .IN4(n2467), 
        .Q(n494) );
  AO22X1 U517 ( .IN1(n2466), .IN2(n2526), .IN3(\regf[14][0] ), .IN4(n2464), 
        .Q(n495) );
  AO22X1 U518 ( .IN1(n2465), .IN2(n2529), .IN3(\regf[14][1] ), .IN4(n2464), 
        .Q(n496) );
  AO22X1 U519 ( .IN1(n2466), .IN2(n2532), .IN3(\regf[14][2] ), .IN4(n2464), 
        .Q(n497) );
  AO22X1 U520 ( .IN1(n2465), .IN2(n2535), .IN3(\regf[14][3] ), .IN4(n2464), 
        .Q(n498) );
  AO22X1 U521 ( .IN1(n2465), .IN2(n2538), .IN3(\regf[14][4] ), .IN4(n2464), 
        .Q(n499) );
  AO22X1 U522 ( .IN1(n2466), .IN2(n2541), .IN3(\regf[14][5] ), .IN4(n2464), 
        .Q(n500) );
  AO22X1 U523 ( .IN1(n2465), .IN2(n2544), .IN3(\regf[14][6] ), .IN4(n2464), 
        .Q(n501) );
  AO22X1 U524 ( .IN1(n2465), .IN2(n2547), .IN3(\regf[14][7] ), .IN4(n2464), 
        .Q(n502) );
  AO22X1 U525 ( .IN1(n2466), .IN2(n2550), .IN3(\regf[14][8] ), .IN4(n2464), 
        .Q(n503) );
  AO22X1 U526 ( .IN1(n2466), .IN2(n2553), .IN3(\regf[14][9] ), .IN4(n2464), 
        .Q(n504) );
  AO22X1 U527 ( .IN1(n2465), .IN2(n2556), .IN3(\regf[14][10] ), .IN4(n2464), 
        .Q(n505) );
  AO22X1 U528 ( .IN1(n2465), .IN2(n2559), .IN3(\regf[14][11] ), .IN4(n2464), 
        .Q(n506) );
  AO22X1 U529 ( .IN1(n2465), .IN2(n2562), .IN3(\regf[14][12] ), .IN4(n2464), 
        .Q(n507) );
  AO22X1 U530 ( .IN1(n2465), .IN2(n2565), .IN3(\regf[14][13] ), .IN4(n2463), 
        .Q(n508) );
  AO22X1 U531 ( .IN1(n2465), .IN2(n2568), .IN3(\regf[14][14] ), .IN4(n59), .Q(
        n509) );
  AO22X1 U532 ( .IN1(n2465), .IN2(n2571), .IN3(\regf[14][15] ), .IN4(n59), .Q(
        n510) );
  AO22X1 U533 ( .IN1(n2465), .IN2(n2574), .IN3(\regf[14][16] ), .IN4(n59), .Q(
        n511) );
  AO22X1 U534 ( .IN1(n2465), .IN2(n2577), .IN3(\regf[14][17] ), .IN4(n59), .Q(
        n512) );
  AO22X1 U535 ( .IN1(n2466), .IN2(n2580), .IN3(\regf[14][18] ), .IN4(n59), .Q(
        n513) );
  AO22X1 U536 ( .IN1(n2465), .IN2(n2583), .IN3(\regf[14][19] ), .IN4(n59), .Q(
        n514) );
  AO22X1 U537 ( .IN1(n2466), .IN2(n2586), .IN3(\regf[14][20] ), .IN4(n2463), 
        .Q(n515) );
  AO22X1 U538 ( .IN1(n2465), .IN2(n2589), .IN3(\regf[14][21] ), .IN4(n2463), 
        .Q(n516) );
  AO22X1 U539 ( .IN1(n2466), .IN2(n2592), .IN3(\regf[14][22] ), .IN4(n2463), 
        .Q(n517) );
  AO22X1 U540 ( .IN1(n2465), .IN2(n2595), .IN3(\regf[14][23] ), .IN4(n2463), 
        .Q(n518) );
  AO22X1 U541 ( .IN1(n2466), .IN2(n2598), .IN3(\regf[14][24] ), .IN4(n2463), 
        .Q(n519) );
  AO22X1 U542 ( .IN1(n2466), .IN2(n2601), .IN3(\regf[14][25] ), .IN4(n2463), 
        .Q(n520) );
  AO22X1 U543 ( .IN1(n2466), .IN2(n2604), .IN3(\regf[14][26] ), .IN4(n2463), 
        .Q(n521) );
  AO22X1 U544 ( .IN1(n2466), .IN2(n2607), .IN3(\regf[14][27] ), .IN4(n2463), 
        .Q(n522) );
  AO22X1 U545 ( .IN1(n2466), .IN2(n2610), .IN3(\regf[14][28] ), .IN4(n2463), 
        .Q(n523) );
  AO22X1 U546 ( .IN1(n2466), .IN2(n2613), .IN3(\regf[14][29] ), .IN4(n2463), 
        .Q(n524) );
  AO22X1 U547 ( .IN1(n2466), .IN2(n2616), .IN3(\regf[14][30] ), .IN4(n2463), 
        .Q(n525) );
  AO22X1 U548 ( .IN1(n2466), .IN2(n2619), .IN3(\regf[14][31] ), .IN4(n2463), 
        .Q(n526) );
  AO22X1 U549 ( .IN1(n2462), .IN2(n2526), .IN3(\regf[15][0] ), .IN4(n2460), 
        .Q(n527) );
  AO22X1 U550 ( .IN1(n2461), .IN2(n2529), .IN3(\regf[15][1] ), .IN4(n2460), 
        .Q(n528) );
  AO22X1 U551 ( .IN1(n2462), .IN2(n2532), .IN3(\regf[15][2] ), .IN4(n2460), 
        .Q(n529) );
  AO22X1 U552 ( .IN1(n2461), .IN2(n2535), .IN3(\regf[15][3] ), .IN4(n2460), 
        .Q(n530) );
  AO22X1 U553 ( .IN1(n2461), .IN2(n2538), .IN3(\regf[15][4] ), .IN4(n2460), 
        .Q(n531) );
  AO22X1 U554 ( .IN1(n2462), .IN2(n2541), .IN3(\regf[15][5] ), .IN4(n2460), 
        .Q(n532) );
  AO22X1 U555 ( .IN1(n2461), .IN2(n2544), .IN3(\regf[15][6] ), .IN4(n2460), 
        .Q(n533) );
  AO22X1 U556 ( .IN1(n2461), .IN2(n2547), .IN3(\regf[15][7] ), .IN4(n2460), 
        .Q(n534) );
  AO22X1 U557 ( .IN1(n2462), .IN2(n2550), .IN3(\regf[15][8] ), .IN4(n2460), 
        .Q(n535) );
  AO22X1 U558 ( .IN1(n2462), .IN2(n2553), .IN3(\regf[15][9] ), .IN4(n2460), 
        .Q(n536) );
  AO22X1 U559 ( .IN1(n2461), .IN2(n2556), .IN3(\regf[15][10] ), .IN4(n2460), 
        .Q(n537) );
  AO22X1 U560 ( .IN1(n2461), .IN2(n2559), .IN3(\regf[15][11] ), .IN4(n2460), 
        .Q(n538) );
  AO22X1 U561 ( .IN1(n2461), .IN2(n2562), .IN3(\regf[15][12] ), .IN4(n2460), 
        .Q(n539) );
  AO22X1 U562 ( .IN1(n2461), .IN2(n2565), .IN3(\regf[15][13] ), .IN4(n2459), 
        .Q(n540) );
  AO22X1 U563 ( .IN1(n2461), .IN2(n2568), .IN3(\regf[15][14] ), .IN4(n60), .Q(
        n541) );
  AO22X1 U564 ( .IN1(n2461), .IN2(n2571), .IN3(\regf[15][15] ), .IN4(n60), .Q(
        n542) );
  AO22X1 U565 ( .IN1(n2461), .IN2(n2574), .IN3(\regf[15][16] ), .IN4(n60), .Q(
        n543) );
  AO22X1 U566 ( .IN1(n2461), .IN2(n2577), .IN3(\regf[15][17] ), .IN4(n60), .Q(
        n544) );
  AO22X1 U567 ( .IN1(n2462), .IN2(n2580), .IN3(\regf[15][18] ), .IN4(n60), .Q(
        n545) );
  AO22X1 U568 ( .IN1(n2461), .IN2(n2583), .IN3(\regf[15][19] ), .IN4(n60), .Q(
        n546) );
  AO22X1 U569 ( .IN1(n2462), .IN2(n2586), .IN3(\regf[15][20] ), .IN4(n2459), 
        .Q(n547) );
  AO22X1 U570 ( .IN1(n2461), .IN2(n2589), .IN3(\regf[15][21] ), .IN4(n2459), 
        .Q(n548) );
  AO22X1 U571 ( .IN1(n2462), .IN2(n2592), .IN3(\regf[15][22] ), .IN4(n2459), 
        .Q(n549) );
  AO22X1 U572 ( .IN1(n2461), .IN2(n2595), .IN3(\regf[15][23] ), .IN4(n2459), 
        .Q(n550) );
  AO22X1 U573 ( .IN1(n2462), .IN2(n2598), .IN3(\regf[15][24] ), .IN4(n2459), 
        .Q(n551) );
  AO22X1 U574 ( .IN1(n2462), .IN2(n2601), .IN3(\regf[15][25] ), .IN4(n2459), 
        .Q(n552) );
  AO22X1 U575 ( .IN1(n2462), .IN2(n2604), .IN3(\regf[15][26] ), .IN4(n2459), 
        .Q(n553) );
  AO22X1 U576 ( .IN1(n2462), .IN2(n2607), .IN3(\regf[15][27] ), .IN4(n2459), 
        .Q(n554) );
  AO22X1 U577 ( .IN1(n2462), .IN2(n2610), .IN3(\regf[15][28] ), .IN4(n2459), 
        .Q(n555) );
  AO22X1 U578 ( .IN1(n2462), .IN2(n2613), .IN3(\regf[15][29] ), .IN4(n2459), 
        .Q(n556) );
  AO22X1 U579 ( .IN1(n2462), .IN2(n2616), .IN3(\regf[15][30] ), .IN4(n2459), 
        .Q(n557) );
  AO22X1 U580 ( .IN1(n2462), .IN2(n2619), .IN3(\regf[15][31] ), .IN4(n2459), 
        .Q(n558) );
  AO22X1 U582 ( .IN1(n2456), .IN2(n2526), .IN3(\regf[16][0] ), .IN4(n61), .Q(
        n559) );
  AO22X1 U583 ( .IN1(n2456), .IN2(n2529), .IN3(\regf[16][1] ), .IN4(n61), .Q(
        n560) );
  AO22X1 U584 ( .IN1(n2456), .IN2(n2532), .IN3(\regf[16][2] ), .IN4(n61), .Q(
        n561) );
  AO22X1 U585 ( .IN1(n2456), .IN2(n2535), .IN3(\regf[16][3] ), .IN4(n61), .Q(
        n562) );
  AO22X1 U586 ( .IN1(n2457), .IN2(n2538), .IN3(\regf[16][4] ), .IN4(n61), .Q(
        n563) );
  AO22X1 U587 ( .IN1(n2458), .IN2(n2541), .IN3(\regf[16][5] ), .IN4(n61), .Q(
        n564) );
  AO22X1 U588 ( .IN1(n2458), .IN2(n2544), .IN3(\regf[16][6] ), .IN4(n61), .Q(
        n565) );
  AO22X1 U589 ( .IN1(n2457), .IN2(n2547), .IN3(\regf[16][7] ), .IN4(n61), .Q(
        n566) );
  AO22X1 U590 ( .IN1(n2458), .IN2(n2550), .IN3(\regf[16][8] ), .IN4(n2455), 
        .Q(n567) );
  AO22X1 U591 ( .IN1(n2458), .IN2(n2553), .IN3(\regf[16][9] ), .IN4(n2455), 
        .Q(n568) );
  AO22X1 U592 ( .IN1(n2457), .IN2(n2556), .IN3(\regf[16][10] ), .IN4(n2455), 
        .Q(n569) );
  AO22X1 U593 ( .IN1(n2457), .IN2(n2559), .IN3(\regf[16][11] ), .IN4(n2455), 
        .Q(n570) );
  AO22X1 U594 ( .IN1(n2457), .IN2(n2562), .IN3(\regf[16][12] ), .IN4(n2455), 
        .Q(n571) );
  AO22X1 U595 ( .IN1(n2457), .IN2(n2565), .IN3(\regf[16][13] ), .IN4(n2455), 
        .Q(n572) );
  AO22X1 U596 ( .IN1(n2457), .IN2(n2568), .IN3(\regf[16][14] ), .IN4(n2455), 
        .Q(n573) );
  AO22X1 U597 ( .IN1(n2457), .IN2(n2571), .IN3(\regf[16][15] ), .IN4(n2455), 
        .Q(n574) );
  AO22X1 U598 ( .IN1(n2457), .IN2(n2574), .IN3(\regf[16][16] ), .IN4(n2455), 
        .Q(n575) );
  AO22X1 U599 ( .IN1(n2457), .IN2(n2577), .IN3(\regf[16][17] ), .IN4(n2455), 
        .Q(n576) );
  AO22X1 U600 ( .IN1(n2457), .IN2(n2580), .IN3(\regf[16][18] ), .IN4(n2455), 
        .Q(n577) );
  AO22X1 U601 ( .IN1(n2458), .IN2(n2583), .IN3(\regf[16][19] ), .IN4(n2455), 
        .Q(n578) );
  AO22X1 U602 ( .IN1(n2457), .IN2(n2586), .IN3(\regf[16][20] ), .IN4(n2454), 
        .Q(n579) );
  AO22X1 U603 ( .IN1(n2458), .IN2(n2589), .IN3(\regf[16][21] ), .IN4(n2454), 
        .Q(n580) );
  AO22X1 U604 ( .IN1(n2457), .IN2(n2592), .IN3(\regf[16][22] ), .IN4(n2454), 
        .Q(n581) );
  AO22X1 U605 ( .IN1(n2458), .IN2(n2595), .IN3(\regf[16][23] ), .IN4(n2454), 
        .Q(n582) );
  AO22X1 U606 ( .IN1(n2457), .IN2(n2598), .IN3(\regf[16][24] ), .IN4(n2454), 
        .Q(n583) );
  AO22X1 U607 ( .IN1(n2458), .IN2(n2601), .IN3(\regf[16][25] ), .IN4(n2454), 
        .Q(n584) );
  AO22X1 U608 ( .IN1(n2458), .IN2(n2604), .IN3(\regf[16][26] ), .IN4(n2454), 
        .Q(n585) );
  AO22X1 U609 ( .IN1(n2458), .IN2(n2607), .IN3(\regf[16][27] ), .IN4(n2454), 
        .Q(n586) );
  AO22X1 U610 ( .IN1(n2458), .IN2(n2610), .IN3(\regf[16][28] ), .IN4(n2454), 
        .Q(n587) );
  AO22X1 U611 ( .IN1(n2458), .IN2(n2613), .IN3(\regf[16][29] ), .IN4(n2454), 
        .Q(n588) );
  AO22X1 U612 ( .IN1(n2458), .IN2(n2616), .IN3(\regf[16][30] ), .IN4(n2454), 
        .Q(n589) );
  AO22X1 U613 ( .IN1(n2458), .IN2(n2619), .IN3(\regf[16][31] ), .IN4(n2454), 
        .Q(n590) );
  AO22X1 U614 ( .IN1(n2451), .IN2(n2526), .IN3(\regf[17][0] ), .IN4(n63), .Q(
        n591) );
  AO22X1 U615 ( .IN1(n2451), .IN2(n2529), .IN3(\regf[17][1] ), .IN4(n63), .Q(
        n592) );
  AO22X1 U616 ( .IN1(n2451), .IN2(n2532), .IN3(\regf[17][2] ), .IN4(n63), .Q(
        n593) );
  AO22X1 U617 ( .IN1(n2451), .IN2(n2535), .IN3(\regf[17][3] ), .IN4(n63), .Q(
        n594) );
  AO22X1 U618 ( .IN1(n2452), .IN2(n2538), .IN3(\regf[17][4] ), .IN4(n63), .Q(
        n595) );
  AO22X1 U619 ( .IN1(n2453), .IN2(n2541), .IN3(\regf[17][5] ), .IN4(n63), .Q(
        n596) );
  AO22X1 U620 ( .IN1(n2453), .IN2(n2544), .IN3(\regf[17][6] ), .IN4(n63), .Q(
        n597) );
  AO22X1 U621 ( .IN1(n2452), .IN2(n2547), .IN3(\regf[17][7] ), .IN4(n63), .Q(
        n598) );
  AO22X1 U622 ( .IN1(n2453), .IN2(n2550), .IN3(\regf[17][8] ), .IN4(n2450), 
        .Q(n599) );
  AO22X1 U623 ( .IN1(n2453), .IN2(n2553), .IN3(\regf[17][9] ), .IN4(n2450), 
        .Q(n600) );
  AO22X1 U624 ( .IN1(n2452), .IN2(n2556), .IN3(\regf[17][10] ), .IN4(n2450), 
        .Q(n601) );
  AO22X1 U625 ( .IN1(n2452), .IN2(n2559), .IN3(\regf[17][11] ), .IN4(n2450), 
        .Q(n602) );
  AO22X1 U626 ( .IN1(n2452), .IN2(n2562), .IN3(\regf[17][12] ), .IN4(n2450), 
        .Q(n603) );
  AO22X1 U627 ( .IN1(n2452), .IN2(n2565), .IN3(\regf[17][13] ), .IN4(n2450), 
        .Q(n604) );
  AO22X1 U628 ( .IN1(n2452), .IN2(n2568), .IN3(\regf[17][14] ), .IN4(n2450), 
        .Q(n605) );
  AO22X1 U629 ( .IN1(n2452), .IN2(n2571), .IN3(\regf[17][15] ), .IN4(n2450), 
        .Q(n606) );
  AO22X1 U630 ( .IN1(n2452), .IN2(n2574), .IN3(\regf[17][16] ), .IN4(n2450), 
        .Q(n607) );
  AO22X1 U631 ( .IN1(n2452), .IN2(n2577), .IN3(\regf[17][17] ), .IN4(n2450), 
        .Q(n608) );
  AO22X1 U632 ( .IN1(n2452), .IN2(n2580), .IN3(\regf[17][18] ), .IN4(n2450), 
        .Q(n609) );
  AO22X1 U633 ( .IN1(n2453), .IN2(n2583), .IN3(\regf[17][19] ), .IN4(n2450), 
        .Q(n610) );
  AO22X1 U634 ( .IN1(n2452), .IN2(n2586), .IN3(\regf[17][20] ), .IN4(n2449), 
        .Q(n611) );
  AO22X1 U635 ( .IN1(n2453), .IN2(n2589), .IN3(\regf[17][21] ), .IN4(n2449), 
        .Q(n612) );
  AO22X1 U636 ( .IN1(n2452), .IN2(n2592), .IN3(\regf[17][22] ), .IN4(n2449), 
        .Q(n613) );
  AO22X1 U637 ( .IN1(n2453), .IN2(n2595), .IN3(\regf[17][23] ), .IN4(n2449), 
        .Q(n614) );
  AO22X1 U638 ( .IN1(n2452), .IN2(n2598), .IN3(\regf[17][24] ), .IN4(n2449), 
        .Q(n615) );
  AO22X1 U639 ( .IN1(n2453), .IN2(n2601), .IN3(\regf[17][25] ), .IN4(n2449), 
        .Q(n616) );
  AO22X1 U640 ( .IN1(n2453), .IN2(n2604), .IN3(\regf[17][26] ), .IN4(n2449), 
        .Q(n617) );
  AO22X1 U641 ( .IN1(n2453), .IN2(n2607), .IN3(\regf[17][27] ), .IN4(n2449), 
        .Q(n618) );
  AO22X1 U642 ( .IN1(n2453), .IN2(n2610), .IN3(\regf[17][28] ), .IN4(n2449), 
        .Q(n619) );
  AO22X1 U643 ( .IN1(n2453), .IN2(n2613), .IN3(\regf[17][29] ), .IN4(n2449), 
        .Q(n620) );
  AO22X1 U644 ( .IN1(n2453), .IN2(n2616), .IN3(\regf[17][30] ), .IN4(n2449), 
        .Q(n621) );
  AO22X1 U645 ( .IN1(n2453), .IN2(n2619), .IN3(\regf[17][31] ), .IN4(n2449), 
        .Q(n622) );
  AO22X1 U646 ( .IN1(n2446), .IN2(n2526), .IN3(\regf[18][0] ), .IN4(n64), .Q(
        n623) );
  AO22X1 U647 ( .IN1(n2446), .IN2(n2529), .IN3(\regf[18][1] ), .IN4(n64), .Q(
        n624) );
  AO22X1 U648 ( .IN1(n2446), .IN2(n2532), .IN3(\regf[18][2] ), .IN4(n64), .Q(
        n625) );
  AO22X1 U649 ( .IN1(n2446), .IN2(n2535), .IN3(\regf[18][3] ), .IN4(n64), .Q(
        n626) );
  AO22X1 U650 ( .IN1(n2447), .IN2(n2538), .IN3(\regf[18][4] ), .IN4(n64), .Q(
        n627) );
  AO22X1 U651 ( .IN1(n2448), .IN2(n2541), .IN3(\regf[18][5] ), .IN4(n64), .Q(
        n628) );
  AO22X1 U652 ( .IN1(n2448), .IN2(n2544), .IN3(\regf[18][6] ), .IN4(n64), .Q(
        n629) );
  AO22X1 U653 ( .IN1(n2447), .IN2(n2547), .IN3(\regf[18][7] ), .IN4(n64), .Q(
        n630) );
  AO22X1 U654 ( .IN1(n2448), .IN2(n2550), .IN3(\regf[18][8] ), .IN4(n2445), 
        .Q(n631) );
  AO22X1 U655 ( .IN1(n2448), .IN2(n2553), .IN3(\regf[18][9] ), .IN4(n2445), 
        .Q(n632) );
  AO22X1 U656 ( .IN1(n2447), .IN2(n2556), .IN3(\regf[18][10] ), .IN4(n2445), 
        .Q(n633) );
  AO22X1 U657 ( .IN1(n2447), .IN2(n2559), .IN3(\regf[18][11] ), .IN4(n2445), 
        .Q(n634) );
  AO22X1 U658 ( .IN1(n2447), .IN2(n2562), .IN3(\regf[18][12] ), .IN4(n2445), 
        .Q(n635) );
  AO22X1 U659 ( .IN1(n2447), .IN2(n2565), .IN3(\regf[18][13] ), .IN4(n2445), 
        .Q(n636) );
  AO22X1 U660 ( .IN1(n2447), .IN2(n2568), .IN3(\regf[18][14] ), .IN4(n2445), 
        .Q(n637) );
  AO22X1 U661 ( .IN1(n2447), .IN2(n2571), .IN3(\regf[18][15] ), .IN4(n2445), 
        .Q(n638) );
  AO22X1 U662 ( .IN1(n2447), .IN2(n2574), .IN3(\regf[18][16] ), .IN4(n2445), 
        .Q(n639) );
  AO22X1 U663 ( .IN1(n2447), .IN2(n2577), .IN3(\regf[18][17] ), .IN4(n2445), 
        .Q(n640) );
  AO22X1 U664 ( .IN1(n2447), .IN2(n2580), .IN3(\regf[18][18] ), .IN4(n2445), 
        .Q(n641) );
  AO22X1 U665 ( .IN1(n2448), .IN2(n2583), .IN3(\regf[18][19] ), .IN4(n2445), 
        .Q(n642) );
  AO22X1 U666 ( .IN1(n2447), .IN2(n2586), .IN3(\regf[18][20] ), .IN4(n2444), 
        .Q(n643) );
  AO22X1 U667 ( .IN1(n2448), .IN2(n2589), .IN3(\regf[18][21] ), .IN4(n2444), 
        .Q(n644) );
  AO22X1 U668 ( .IN1(n2447), .IN2(n2592), .IN3(\regf[18][22] ), .IN4(n2444), 
        .Q(n645) );
  AO22X1 U669 ( .IN1(n2448), .IN2(n2595), .IN3(\regf[18][23] ), .IN4(n2444), 
        .Q(n646) );
  AO22X1 U670 ( .IN1(n2447), .IN2(n2598), .IN3(\regf[18][24] ), .IN4(n2444), 
        .Q(n647) );
  AO22X1 U671 ( .IN1(n2448), .IN2(n2601), .IN3(\regf[18][25] ), .IN4(n2444), 
        .Q(n648) );
  AO22X1 U672 ( .IN1(n2448), .IN2(n2604), .IN3(\regf[18][26] ), .IN4(n2444), 
        .Q(n649) );
  AO22X1 U673 ( .IN1(n2448), .IN2(n2607), .IN3(\regf[18][27] ), .IN4(n2444), 
        .Q(n650) );
  AO22X1 U674 ( .IN1(n2448), .IN2(n2610), .IN3(\regf[18][28] ), .IN4(n2444), 
        .Q(n651) );
  AO22X1 U675 ( .IN1(n2448), .IN2(n2613), .IN3(\regf[18][29] ), .IN4(n2444), 
        .Q(n652) );
  AO22X1 U676 ( .IN1(n2448), .IN2(n2616), .IN3(\regf[18][30] ), .IN4(n2444), 
        .Q(n653) );
  AO22X1 U677 ( .IN1(n2448), .IN2(n2619), .IN3(\regf[18][31] ), .IN4(n2444), 
        .Q(n654) );
  AO22X1 U678 ( .IN1(n2441), .IN2(n2526), .IN3(\regf[19][0] ), .IN4(n65), .Q(
        n655) );
  AO22X1 U679 ( .IN1(n2441), .IN2(n2529), .IN3(\regf[19][1] ), .IN4(n65), .Q(
        n656) );
  AO22X1 U680 ( .IN1(n2441), .IN2(n2532), .IN3(\regf[19][2] ), .IN4(n65), .Q(
        n657) );
  AO22X1 U681 ( .IN1(n2441), .IN2(n2535), .IN3(\regf[19][3] ), .IN4(n65), .Q(
        n658) );
  AO22X1 U682 ( .IN1(n2442), .IN2(n2538), .IN3(\regf[19][4] ), .IN4(n65), .Q(
        n659) );
  AO22X1 U683 ( .IN1(n2443), .IN2(n2541), .IN3(\regf[19][5] ), .IN4(n65), .Q(
        n660) );
  AO22X1 U684 ( .IN1(n2443), .IN2(n2544), .IN3(\regf[19][6] ), .IN4(n65), .Q(
        n661) );
  AO22X1 U685 ( .IN1(n2442), .IN2(n2547), .IN3(\regf[19][7] ), .IN4(n65), .Q(
        n662) );
  AO22X1 U686 ( .IN1(n2443), .IN2(n2550), .IN3(\regf[19][8] ), .IN4(n2440), 
        .Q(n663) );
  AO22X1 U687 ( .IN1(n2443), .IN2(n2553), .IN3(\regf[19][9] ), .IN4(n2440), 
        .Q(n664) );
  AO22X1 U688 ( .IN1(n2442), .IN2(n2556), .IN3(\regf[19][10] ), .IN4(n2440), 
        .Q(n665) );
  AO22X1 U689 ( .IN1(n2442), .IN2(n2559), .IN3(\regf[19][11] ), .IN4(n2440), 
        .Q(n666) );
  AO22X1 U690 ( .IN1(n2442), .IN2(n2562), .IN3(\regf[19][12] ), .IN4(n2440), 
        .Q(n667) );
  AO22X1 U691 ( .IN1(n2442), .IN2(n2565), .IN3(\regf[19][13] ), .IN4(n2440), 
        .Q(n668) );
  AO22X1 U692 ( .IN1(n2442), .IN2(n2568), .IN3(\regf[19][14] ), .IN4(n2440), 
        .Q(n669) );
  AO22X1 U693 ( .IN1(n2442), .IN2(n2571), .IN3(\regf[19][15] ), .IN4(n2440), 
        .Q(n670) );
  AO22X1 U694 ( .IN1(n2442), .IN2(n2574), .IN3(\regf[19][16] ), .IN4(n2440), 
        .Q(n671) );
  AO22X1 U695 ( .IN1(n2442), .IN2(n2577), .IN3(\regf[19][17] ), .IN4(n2440), 
        .Q(n672) );
  AO22X1 U696 ( .IN1(n2442), .IN2(n2580), .IN3(\regf[19][18] ), .IN4(n2440), 
        .Q(n673) );
  AO22X1 U697 ( .IN1(n2443), .IN2(n2583), .IN3(\regf[19][19] ), .IN4(n2440), 
        .Q(n674) );
  AO22X1 U698 ( .IN1(n2442), .IN2(n2586), .IN3(\regf[19][20] ), .IN4(n2439), 
        .Q(n675) );
  AO22X1 U699 ( .IN1(n2443), .IN2(n2589), .IN3(\regf[19][21] ), .IN4(n2439), 
        .Q(n676) );
  AO22X1 U700 ( .IN1(n2442), .IN2(n2592), .IN3(\regf[19][22] ), .IN4(n2439), 
        .Q(n677) );
  AO22X1 U701 ( .IN1(n2443), .IN2(n2595), .IN3(\regf[19][23] ), .IN4(n2439), 
        .Q(n678) );
  AO22X1 U702 ( .IN1(n2442), .IN2(n2598), .IN3(\regf[19][24] ), .IN4(n2439), 
        .Q(n679) );
  AO22X1 U703 ( .IN1(n2443), .IN2(n2601), .IN3(\regf[19][25] ), .IN4(n2439), 
        .Q(n680) );
  AO22X1 U704 ( .IN1(n2443), .IN2(n2604), .IN3(\regf[19][26] ), .IN4(n2439), 
        .Q(n681) );
  AO22X1 U705 ( .IN1(n2443), .IN2(n2607), .IN3(\regf[19][27] ), .IN4(n2439), 
        .Q(n682) );
  AO22X1 U706 ( .IN1(n2443), .IN2(n2610), .IN3(\regf[19][28] ), .IN4(n2439), 
        .Q(n683) );
  AO22X1 U707 ( .IN1(n2443), .IN2(n2613), .IN3(\regf[19][29] ), .IN4(n2439), 
        .Q(n684) );
  AO22X1 U708 ( .IN1(n2443), .IN2(n2616), .IN3(\regf[19][30] ), .IN4(n2439), 
        .Q(n685) );
  AO22X1 U709 ( .IN1(n2443), .IN2(n2619), .IN3(\regf[19][31] ), .IN4(n2439), 
        .Q(n686) );
  AO22X1 U710 ( .IN1(n2436), .IN2(n2526), .IN3(\regf[20][0] ), .IN4(n66), .Q(
        n687) );
  AO22X1 U711 ( .IN1(n2436), .IN2(n2529), .IN3(\regf[20][1] ), .IN4(n66), .Q(
        n688) );
  AO22X1 U712 ( .IN1(n2436), .IN2(n2532), .IN3(\regf[20][2] ), .IN4(n66), .Q(
        n689) );
  AO22X1 U713 ( .IN1(n2436), .IN2(n2535), .IN3(\regf[20][3] ), .IN4(n66), .Q(
        n690) );
  AO22X1 U714 ( .IN1(n2437), .IN2(n2538), .IN3(\regf[20][4] ), .IN4(n66), .Q(
        n691) );
  AO22X1 U715 ( .IN1(n2438), .IN2(n2541), .IN3(\regf[20][5] ), .IN4(n66), .Q(
        n692) );
  AO22X1 U716 ( .IN1(n2438), .IN2(n2544), .IN3(\regf[20][6] ), .IN4(n66), .Q(
        n693) );
  AO22X1 U717 ( .IN1(n2437), .IN2(n2547), .IN3(\regf[20][7] ), .IN4(n66), .Q(
        n694) );
  AO22X1 U718 ( .IN1(n2438), .IN2(n2550), .IN3(\regf[20][8] ), .IN4(n2435), 
        .Q(n695) );
  AO22X1 U719 ( .IN1(n2438), .IN2(n2553), .IN3(\regf[20][9] ), .IN4(n2435), 
        .Q(n696) );
  AO22X1 U720 ( .IN1(n2437), .IN2(n2556), .IN3(\regf[20][10] ), .IN4(n2435), 
        .Q(n697) );
  AO22X1 U721 ( .IN1(n2437), .IN2(n2559), .IN3(\regf[20][11] ), .IN4(n2435), 
        .Q(n698) );
  AO22X1 U722 ( .IN1(n2437), .IN2(n2562), .IN3(\regf[20][12] ), .IN4(n2435), 
        .Q(n699) );
  AO22X1 U723 ( .IN1(n2437), .IN2(n2565), .IN3(\regf[20][13] ), .IN4(n2435), 
        .Q(n700) );
  AO22X1 U724 ( .IN1(n2437), .IN2(n2568), .IN3(\regf[20][14] ), .IN4(n2435), 
        .Q(n701) );
  AO22X1 U725 ( .IN1(n2437), .IN2(n2571), .IN3(\regf[20][15] ), .IN4(n2435), 
        .Q(n702) );
  AO22X1 U726 ( .IN1(n2437), .IN2(n2574), .IN3(\regf[20][16] ), .IN4(n2435), 
        .Q(n703) );
  AO22X1 U727 ( .IN1(n2437), .IN2(n2577), .IN3(\regf[20][17] ), .IN4(n2435), 
        .Q(n704) );
  AO22X1 U728 ( .IN1(n2437), .IN2(n2580), .IN3(\regf[20][18] ), .IN4(n2435), 
        .Q(n705) );
  AO22X1 U729 ( .IN1(n2438), .IN2(n2583), .IN3(\regf[20][19] ), .IN4(n2435), 
        .Q(n706) );
  AO22X1 U730 ( .IN1(n2437), .IN2(n2586), .IN3(\regf[20][20] ), .IN4(n2434), 
        .Q(n707) );
  AO22X1 U731 ( .IN1(n2438), .IN2(n2589), .IN3(\regf[20][21] ), .IN4(n2434), 
        .Q(n708) );
  AO22X1 U732 ( .IN1(n2437), .IN2(n2592), .IN3(\regf[20][22] ), .IN4(n2434), 
        .Q(n709) );
  AO22X1 U733 ( .IN1(n2438), .IN2(n2595), .IN3(\regf[20][23] ), .IN4(n2434), 
        .Q(n710) );
  AO22X1 U734 ( .IN1(n2437), .IN2(n2598), .IN3(\regf[20][24] ), .IN4(n2434), 
        .Q(n711) );
  AO22X1 U735 ( .IN1(n2438), .IN2(n2601), .IN3(\regf[20][25] ), .IN4(n2434), 
        .Q(n712) );
  AO22X1 U736 ( .IN1(n2438), .IN2(n2604), .IN3(\regf[20][26] ), .IN4(n2434), 
        .Q(n713) );
  AO22X1 U737 ( .IN1(n2438), .IN2(n2607), .IN3(\regf[20][27] ), .IN4(n2434), 
        .Q(n714) );
  AO22X1 U738 ( .IN1(n2438), .IN2(n2610), .IN3(\regf[20][28] ), .IN4(n2434), 
        .Q(n715) );
  AO22X1 U739 ( .IN1(n2438), .IN2(n2613), .IN3(\regf[20][29] ), .IN4(n2434), 
        .Q(n716) );
  AO22X1 U740 ( .IN1(n2438), .IN2(n2616), .IN3(\regf[20][30] ), .IN4(n2434), 
        .Q(n717) );
  AO22X1 U741 ( .IN1(n2438), .IN2(n2619), .IN3(\regf[20][31] ), .IN4(n2434), 
        .Q(n718) );
  AO22X1 U742 ( .IN1(n2431), .IN2(n2526), .IN3(\regf[21][0] ), .IN4(n67), .Q(
        n719) );
  AO22X1 U743 ( .IN1(n2431), .IN2(n2529), .IN3(\regf[21][1] ), .IN4(n67), .Q(
        n720) );
  AO22X1 U744 ( .IN1(n2431), .IN2(n2532), .IN3(\regf[21][2] ), .IN4(n67), .Q(
        n721) );
  AO22X1 U745 ( .IN1(n2431), .IN2(n2535), .IN3(\regf[21][3] ), .IN4(n67), .Q(
        n722) );
  AO22X1 U746 ( .IN1(n2432), .IN2(n2538), .IN3(\regf[21][4] ), .IN4(n67), .Q(
        n723) );
  AO22X1 U747 ( .IN1(n2433), .IN2(n2541), .IN3(\regf[21][5] ), .IN4(n67), .Q(
        n724) );
  AO22X1 U748 ( .IN1(n2433), .IN2(n2544), .IN3(\regf[21][6] ), .IN4(n67), .Q(
        n725) );
  AO22X1 U749 ( .IN1(n2432), .IN2(n2547), .IN3(\regf[21][7] ), .IN4(n67), .Q(
        n726) );
  AO22X1 U750 ( .IN1(n2433), .IN2(n2550), .IN3(\regf[21][8] ), .IN4(n2430), 
        .Q(n727) );
  AO22X1 U751 ( .IN1(n2433), .IN2(n2553), .IN3(\regf[21][9] ), .IN4(n2430), 
        .Q(n728) );
  AO22X1 U752 ( .IN1(n2432), .IN2(n2556), .IN3(\regf[21][10] ), .IN4(n2430), 
        .Q(n729) );
  AO22X1 U753 ( .IN1(n2432), .IN2(n2559), .IN3(\regf[21][11] ), .IN4(n2430), 
        .Q(n730) );
  AO22X1 U754 ( .IN1(n2432), .IN2(n2562), .IN3(\regf[21][12] ), .IN4(n2430), 
        .Q(n731) );
  AO22X1 U755 ( .IN1(n2432), .IN2(n2565), .IN3(\regf[21][13] ), .IN4(n2430), 
        .Q(n732) );
  AO22X1 U756 ( .IN1(n2432), .IN2(n2568), .IN3(\regf[21][14] ), .IN4(n2430), 
        .Q(n733) );
  AO22X1 U757 ( .IN1(n2432), .IN2(n2571), .IN3(\regf[21][15] ), .IN4(n2430), 
        .Q(n734) );
  AO22X1 U758 ( .IN1(n2432), .IN2(n2574), .IN3(\regf[21][16] ), .IN4(n2430), 
        .Q(n735) );
  AO22X1 U759 ( .IN1(n2432), .IN2(n2577), .IN3(\regf[21][17] ), .IN4(n2430), 
        .Q(n736) );
  AO22X1 U760 ( .IN1(n2432), .IN2(n2580), .IN3(\regf[21][18] ), .IN4(n2430), 
        .Q(n737) );
  AO22X1 U761 ( .IN1(n2433), .IN2(n2583), .IN3(\regf[21][19] ), .IN4(n2430), 
        .Q(n738) );
  AO22X1 U762 ( .IN1(n2432), .IN2(n2586), .IN3(\regf[21][20] ), .IN4(n2429), 
        .Q(n739) );
  AO22X1 U763 ( .IN1(n2433), .IN2(n2589), .IN3(\regf[21][21] ), .IN4(n2429), 
        .Q(n740) );
  AO22X1 U764 ( .IN1(n2432), .IN2(n2592), .IN3(\regf[21][22] ), .IN4(n2429), 
        .Q(n741) );
  AO22X1 U765 ( .IN1(n2433), .IN2(n2595), .IN3(\regf[21][23] ), .IN4(n2429), 
        .Q(n742) );
  AO22X1 U766 ( .IN1(n2432), .IN2(n2598), .IN3(\regf[21][24] ), .IN4(n2429), 
        .Q(n743) );
  AO22X1 U767 ( .IN1(n2433), .IN2(n2601), .IN3(\regf[21][25] ), .IN4(n2429), 
        .Q(n744) );
  AO22X1 U768 ( .IN1(n2433), .IN2(n2604), .IN3(\regf[21][26] ), .IN4(n2429), 
        .Q(n745) );
  AO22X1 U769 ( .IN1(n2433), .IN2(n2607), .IN3(\regf[21][27] ), .IN4(n2429), 
        .Q(n746) );
  AO22X1 U770 ( .IN1(n2433), .IN2(n2610), .IN3(\regf[21][28] ), .IN4(n2429), 
        .Q(n747) );
  AO22X1 U771 ( .IN1(n2433), .IN2(n2613), .IN3(\regf[21][29] ), .IN4(n2429), 
        .Q(n748) );
  AO22X1 U772 ( .IN1(n2433), .IN2(n2616), .IN3(\regf[21][30] ), .IN4(n2429), 
        .Q(n749) );
  AO22X1 U773 ( .IN1(n2433), .IN2(n2619), .IN3(\regf[21][31] ), .IN4(n2429), 
        .Q(n750) );
  AO22X1 U774 ( .IN1(n2426), .IN2(n2526), .IN3(\regf[22][0] ), .IN4(n68), .Q(
        n751) );
  AO22X1 U775 ( .IN1(n2426), .IN2(n2529), .IN3(\regf[22][1] ), .IN4(n68), .Q(
        n752) );
  AO22X1 U776 ( .IN1(n2426), .IN2(n2532), .IN3(\regf[22][2] ), .IN4(n68), .Q(
        n753) );
  AO22X1 U777 ( .IN1(n2426), .IN2(n2535), .IN3(\regf[22][3] ), .IN4(n68), .Q(
        n754) );
  AO22X1 U778 ( .IN1(n2427), .IN2(n2538), .IN3(\regf[22][4] ), .IN4(n68), .Q(
        n755) );
  AO22X1 U779 ( .IN1(n2428), .IN2(n2541), .IN3(\regf[22][5] ), .IN4(n68), .Q(
        n756) );
  AO22X1 U780 ( .IN1(n2428), .IN2(n2544), .IN3(\regf[22][6] ), .IN4(n68), .Q(
        n757) );
  AO22X1 U781 ( .IN1(n2427), .IN2(n2547), .IN3(\regf[22][7] ), .IN4(n68), .Q(
        n758) );
  AO22X1 U782 ( .IN1(n2428), .IN2(n2550), .IN3(\regf[22][8] ), .IN4(n2425), 
        .Q(n759) );
  AO22X1 U783 ( .IN1(n2428), .IN2(n2553), .IN3(\regf[22][9] ), .IN4(n2425), 
        .Q(n760) );
  AO22X1 U784 ( .IN1(n2427), .IN2(n2556), .IN3(\regf[22][10] ), .IN4(n2425), 
        .Q(n761) );
  AO22X1 U785 ( .IN1(n2427), .IN2(n2559), .IN3(\regf[22][11] ), .IN4(n2425), 
        .Q(n762) );
  AO22X1 U786 ( .IN1(n2427), .IN2(n2562), .IN3(\regf[22][12] ), .IN4(n2425), 
        .Q(n763) );
  AO22X1 U787 ( .IN1(n2427), .IN2(n2565), .IN3(\regf[22][13] ), .IN4(n2425), 
        .Q(n764) );
  AO22X1 U788 ( .IN1(n2427), .IN2(n2568), .IN3(\regf[22][14] ), .IN4(n2425), 
        .Q(n765) );
  AO22X1 U789 ( .IN1(n2427), .IN2(n2571), .IN3(\regf[22][15] ), .IN4(n2425), 
        .Q(n766) );
  AO22X1 U790 ( .IN1(n2427), .IN2(n2574), .IN3(\regf[22][16] ), .IN4(n2425), 
        .Q(n767) );
  AO22X1 U791 ( .IN1(n2427), .IN2(n2577), .IN3(\regf[22][17] ), .IN4(n2425), 
        .Q(n768) );
  AO22X1 U792 ( .IN1(n2427), .IN2(n2580), .IN3(\regf[22][18] ), .IN4(n2425), 
        .Q(n769) );
  AO22X1 U793 ( .IN1(n2428), .IN2(n2583), .IN3(\regf[22][19] ), .IN4(n2425), 
        .Q(n770) );
  AO22X1 U794 ( .IN1(n2427), .IN2(n2586), .IN3(\regf[22][20] ), .IN4(n2424), 
        .Q(n771) );
  AO22X1 U795 ( .IN1(n2428), .IN2(n2589), .IN3(\regf[22][21] ), .IN4(n2424), 
        .Q(n772) );
  AO22X1 U796 ( .IN1(n2427), .IN2(n2592), .IN3(\regf[22][22] ), .IN4(n2424), 
        .Q(n773) );
  AO22X1 U797 ( .IN1(n2428), .IN2(n2595), .IN3(\regf[22][23] ), .IN4(n2424), 
        .Q(n774) );
  AO22X1 U798 ( .IN1(n2427), .IN2(n2598), .IN3(\regf[22][24] ), .IN4(n2424), 
        .Q(n775) );
  AO22X1 U799 ( .IN1(n2428), .IN2(n2601), .IN3(\regf[22][25] ), .IN4(n2424), 
        .Q(n776) );
  AO22X1 U800 ( .IN1(n2428), .IN2(n2604), .IN3(\regf[22][26] ), .IN4(n2424), 
        .Q(n777) );
  AO22X1 U801 ( .IN1(n2428), .IN2(n2607), .IN3(\regf[22][27] ), .IN4(n2424), 
        .Q(n778) );
  AO22X1 U802 ( .IN1(n2428), .IN2(n2610), .IN3(\regf[22][28] ), .IN4(n2424), 
        .Q(n779) );
  AO22X1 U803 ( .IN1(n2428), .IN2(n2613), .IN3(\regf[22][29] ), .IN4(n2424), 
        .Q(n780) );
  AO22X1 U804 ( .IN1(n2428), .IN2(n2616), .IN3(\regf[22][30] ), .IN4(n2424), 
        .Q(n781) );
  AO22X1 U805 ( .IN1(n2428), .IN2(n2619), .IN3(\regf[22][31] ), .IN4(n2424), 
        .Q(n782) );
  AO22X1 U806 ( .IN1(n2421), .IN2(n2526), .IN3(\regf[23][0] ), .IN4(n69), .Q(
        n783) );
  AO22X1 U807 ( .IN1(n2421), .IN2(n2529), .IN3(\regf[23][1] ), .IN4(n69), .Q(
        n784) );
  AO22X1 U808 ( .IN1(n2421), .IN2(n2532), .IN3(\regf[23][2] ), .IN4(n69), .Q(
        n785) );
  AO22X1 U809 ( .IN1(n2421), .IN2(n2535), .IN3(\regf[23][3] ), .IN4(n69), .Q(
        n786) );
  AO22X1 U810 ( .IN1(n2422), .IN2(n2538), .IN3(\regf[23][4] ), .IN4(n69), .Q(
        n787) );
  AO22X1 U811 ( .IN1(n2423), .IN2(n2541), .IN3(\regf[23][5] ), .IN4(n69), .Q(
        n788) );
  AO22X1 U812 ( .IN1(n2423), .IN2(n2544), .IN3(\regf[23][6] ), .IN4(n69), .Q(
        n789) );
  AO22X1 U813 ( .IN1(n2422), .IN2(n2547), .IN3(\regf[23][7] ), .IN4(n69), .Q(
        n790) );
  AO22X1 U814 ( .IN1(n2423), .IN2(n2550), .IN3(\regf[23][8] ), .IN4(n2420), 
        .Q(n791) );
  AO22X1 U815 ( .IN1(n2423), .IN2(n2553), .IN3(\regf[23][9] ), .IN4(n2420), 
        .Q(n792) );
  AO22X1 U816 ( .IN1(n2422), .IN2(n2556), .IN3(\regf[23][10] ), .IN4(n2420), 
        .Q(n793) );
  AO22X1 U817 ( .IN1(n2422), .IN2(n2559), .IN3(\regf[23][11] ), .IN4(n2420), 
        .Q(n794) );
  AO22X1 U818 ( .IN1(n2422), .IN2(n2562), .IN3(\regf[23][12] ), .IN4(n2420), 
        .Q(n795) );
  AO22X1 U819 ( .IN1(n2422), .IN2(n2565), .IN3(\regf[23][13] ), .IN4(n2420), 
        .Q(n796) );
  AO22X1 U820 ( .IN1(n2422), .IN2(n2568), .IN3(\regf[23][14] ), .IN4(n2420), 
        .Q(n797) );
  AO22X1 U821 ( .IN1(n2422), .IN2(n2571), .IN3(\regf[23][15] ), .IN4(n2420), 
        .Q(n798) );
  AO22X1 U822 ( .IN1(n2422), .IN2(n2574), .IN3(\regf[23][16] ), .IN4(n2420), 
        .Q(n799) );
  AO22X1 U823 ( .IN1(n2422), .IN2(n2577), .IN3(\regf[23][17] ), .IN4(n2420), 
        .Q(n800) );
  AO22X1 U824 ( .IN1(n2422), .IN2(n2580), .IN3(\regf[23][18] ), .IN4(n2420), 
        .Q(n801) );
  AO22X1 U825 ( .IN1(n2423), .IN2(n2583), .IN3(\regf[23][19] ), .IN4(n2420), 
        .Q(n802) );
  AO22X1 U826 ( .IN1(n2422), .IN2(n2586), .IN3(\regf[23][20] ), .IN4(n2419), 
        .Q(n803) );
  AO22X1 U827 ( .IN1(n2423), .IN2(n2589), .IN3(\regf[23][21] ), .IN4(n2419), 
        .Q(n804) );
  AO22X1 U828 ( .IN1(n2422), .IN2(n2592), .IN3(\regf[23][22] ), .IN4(n2419), 
        .Q(n805) );
  AO22X1 U829 ( .IN1(n2423), .IN2(n2595), .IN3(\regf[23][23] ), .IN4(n2419), 
        .Q(n806) );
  AO22X1 U830 ( .IN1(n2422), .IN2(n2598), .IN3(\regf[23][24] ), .IN4(n2419), 
        .Q(n807) );
  AO22X1 U831 ( .IN1(n2423), .IN2(n2601), .IN3(\regf[23][25] ), .IN4(n2419), 
        .Q(n808) );
  AO22X1 U832 ( .IN1(n2423), .IN2(n2604), .IN3(\regf[23][26] ), .IN4(n2419), 
        .Q(n809) );
  AO22X1 U833 ( .IN1(n2423), .IN2(n2607), .IN3(\regf[23][27] ), .IN4(n2419), 
        .Q(n810) );
  AO22X1 U834 ( .IN1(n2423), .IN2(n2610), .IN3(\regf[23][28] ), .IN4(n2419), 
        .Q(n811) );
  AO22X1 U835 ( .IN1(n2423), .IN2(n2613), .IN3(\regf[23][29] ), .IN4(n2419), 
        .Q(n812) );
  AO22X1 U836 ( .IN1(n2423), .IN2(n2616), .IN3(\regf[23][30] ), .IN4(n2419), 
        .Q(n813) );
  AO22X1 U837 ( .IN1(n2423), .IN2(n2619), .IN3(\regf[23][31] ), .IN4(n2419), 
        .Q(n814) );
  AND3X1 U838 ( .IN1(wr_en), .IN2(n2712), .IN3(wr_addr[4]), .Q(n62) );
  AO22X1 U839 ( .IN1(n2418), .IN2(n2526), .IN3(\regf[24][0] ), .IN4(n2416), 
        .Q(n815) );
  AO22X1 U840 ( .IN1(n2417), .IN2(n2529), .IN3(\regf[24][1] ), .IN4(n2416), 
        .Q(n816) );
  AO22X1 U841 ( .IN1(n2418), .IN2(n2532), .IN3(\regf[24][2] ), .IN4(n2416), 
        .Q(n817) );
  AO22X1 U842 ( .IN1(n2417), .IN2(n2535), .IN3(\regf[24][3] ), .IN4(n2416), 
        .Q(n818) );
  AO22X1 U843 ( .IN1(n2418), .IN2(n2538), .IN3(\regf[24][4] ), .IN4(n2416), 
        .Q(n819) );
  AO22X1 U844 ( .IN1(n2417), .IN2(n2541), .IN3(\regf[24][5] ), .IN4(n2416), 
        .Q(n820) );
  AO22X1 U845 ( .IN1(n2417), .IN2(n2544), .IN3(\regf[24][6] ), .IN4(n2416), 
        .Q(n821) );
  AO22X1 U846 ( .IN1(n2418), .IN2(n2547), .IN3(\regf[24][7] ), .IN4(n2416), 
        .Q(n822) );
  AO22X1 U847 ( .IN1(n2417), .IN2(n2550), .IN3(\regf[24][8] ), .IN4(n2416), 
        .Q(n823) );
  AO22X1 U848 ( .IN1(n2417), .IN2(n2553), .IN3(\regf[24][9] ), .IN4(n2416), 
        .Q(n824) );
  AO22X1 U849 ( .IN1(n2418), .IN2(n2556), .IN3(\regf[24][10] ), .IN4(n2416), 
        .Q(n825) );
  AO22X1 U850 ( .IN1(n2418), .IN2(n2559), .IN3(\regf[24][11] ), .IN4(n2416), 
        .Q(n826) );
  AO22X1 U851 ( .IN1(n2417), .IN2(n2562), .IN3(\regf[24][12] ), .IN4(n2416), 
        .Q(n827) );
  AO22X1 U852 ( .IN1(n2418), .IN2(n2565), .IN3(\regf[24][13] ), .IN4(n2415), 
        .Q(n828) );
  AO22X1 U853 ( .IN1(n2417), .IN2(n2568), .IN3(\regf[24][14] ), .IN4(n70), .Q(
        n829) );
  AO22X1 U854 ( .IN1(n2418), .IN2(n2571), .IN3(\regf[24][15] ), .IN4(n70), .Q(
        n830) );
  AO22X1 U855 ( .IN1(n2417), .IN2(n2574), .IN3(\regf[24][16] ), .IN4(n70), .Q(
        n831) );
  AO22X1 U856 ( .IN1(n2418), .IN2(n2577), .IN3(\regf[24][17] ), .IN4(n70), .Q(
        n832) );
  AO22X1 U857 ( .IN1(n2417), .IN2(n2580), .IN3(\regf[24][18] ), .IN4(n70), .Q(
        n833) );
  AO22X1 U858 ( .IN1(n2417), .IN2(n2583), .IN3(\regf[24][19] ), .IN4(n70), .Q(
        n834) );
  AO22X1 U859 ( .IN1(n2417), .IN2(n2586), .IN3(\regf[24][20] ), .IN4(n2415), 
        .Q(n835) );
  AO22X1 U860 ( .IN1(n2417), .IN2(n2589), .IN3(\regf[24][21] ), .IN4(n2415), 
        .Q(n836) );
  AO22X1 U861 ( .IN1(n2417), .IN2(n2592), .IN3(\regf[24][22] ), .IN4(n2415), 
        .Q(n837) );
  AO22X1 U862 ( .IN1(n2417), .IN2(n2595), .IN3(\regf[24][23] ), .IN4(n2415), 
        .Q(n838) );
  AO22X1 U863 ( .IN1(n2417), .IN2(n2598), .IN3(\regf[24][24] ), .IN4(n2415), 
        .Q(n839) );
  AO22X1 U864 ( .IN1(n2418), .IN2(n2601), .IN3(\regf[24][25] ), .IN4(n2415), 
        .Q(n840) );
  AO22X1 U865 ( .IN1(n2418), .IN2(n2604), .IN3(\regf[24][26] ), .IN4(n2415), 
        .Q(n841) );
  AO22X1 U866 ( .IN1(n2418), .IN2(n2607), .IN3(\regf[24][27] ), .IN4(n2415), 
        .Q(n842) );
  AO22X1 U867 ( .IN1(n2418), .IN2(n2610), .IN3(\regf[24][28] ), .IN4(n2415), 
        .Q(n843) );
  AO22X1 U868 ( .IN1(n2418), .IN2(n2613), .IN3(\regf[24][29] ), .IN4(n2415), 
        .Q(n844) );
  AO22X1 U869 ( .IN1(n2418), .IN2(n2616), .IN3(\regf[24][30] ), .IN4(n2415), 
        .Q(n845) );
  AO22X1 U870 ( .IN1(n2418), .IN2(n2619), .IN3(\regf[24][31] ), .IN4(n2415), 
        .Q(n846) );
  NOR3X0 U871 ( .IN1(wr_addr[1]), .IN2(wr_addr[2]), .IN3(wr_addr[0]), .QN(n36)
         );
  AO22X1 U872 ( .IN1(n2412), .IN2(n2527), .IN3(\regf[25][0] ), .IN4(n2411), 
        .Q(n847) );
  AO22X1 U873 ( .IN1(n2412), .IN2(n2530), .IN3(\regf[25][1] ), .IN4(n2411), 
        .Q(n848) );
  AO22X1 U874 ( .IN1(n2412), .IN2(n2533), .IN3(\regf[25][2] ), .IN4(n2411), 
        .Q(n849) );
  AO22X1 U875 ( .IN1(n2412), .IN2(n2536), .IN3(\regf[25][3] ), .IN4(n2411), 
        .Q(n850) );
  AO22X1 U876 ( .IN1(n2413), .IN2(n2539), .IN3(\regf[25][4] ), .IN4(n2411), 
        .Q(n851) );
  AO22X1 U877 ( .IN1(n2414), .IN2(n2542), .IN3(\regf[25][5] ), .IN4(n2411), 
        .Q(n852) );
  AO22X1 U878 ( .IN1(n2413), .IN2(n2545), .IN3(\regf[25][6] ), .IN4(n2411), 
        .Q(n853) );
  AO22X1 U879 ( .IN1(n2413), .IN2(n2548), .IN3(\regf[25][7] ), .IN4(n2411), 
        .Q(n854) );
  AO22X1 U880 ( .IN1(n2414), .IN2(n2551), .IN3(\regf[25][8] ), .IN4(n2411), 
        .Q(n855) );
  AO22X1 U881 ( .IN1(n2414), .IN2(n2554), .IN3(\regf[25][9] ), .IN4(n2411), 
        .Q(n856) );
  AO22X1 U882 ( .IN1(n2413), .IN2(n2557), .IN3(\regf[25][10] ), .IN4(n2411), 
        .Q(n857) );
  AO22X1 U883 ( .IN1(n2413), .IN2(n2560), .IN3(\regf[25][11] ), .IN4(n2411), 
        .Q(n858) );
  AO22X1 U884 ( .IN1(n2413), .IN2(n2563), .IN3(\regf[25][12] ), .IN4(n2411), 
        .Q(n859) );
  AO22X1 U885 ( .IN1(n2413), .IN2(n2566), .IN3(\regf[25][13] ), .IN4(n2410), 
        .Q(n860) );
  AO22X1 U886 ( .IN1(n2413), .IN2(n2569), .IN3(\regf[25][14] ), .IN4(n72), .Q(
        n861) );
  AO22X1 U887 ( .IN1(n2413), .IN2(n2572), .IN3(\regf[25][15] ), .IN4(n72), .Q(
        n862) );
  AO22X1 U888 ( .IN1(n2413), .IN2(n2575), .IN3(\regf[25][16] ), .IN4(n72), .Q(
        n863) );
  AO22X1 U889 ( .IN1(n2413), .IN2(n2578), .IN3(\regf[25][17] ), .IN4(n72), .Q(
        n864) );
  AO22X1 U890 ( .IN1(n2414), .IN2(n2581), .IN3(\regf[25][18] ), .IN4(n72), .Q(
        n865) );
  AO22X1 U891 ( .IN1(n2413), .IN2(n2584), .IN3(\regf[25][19] ), .IN4(n72), .Q(
        n866) );
  AO22X1 U892 ( .IN1(n2414), .IN2(n2587), .IN3(\regf[25][20] ), .IN4(n2410), 
        .Q(n867) );
  AO22X1 U893 ( .IN1(n2413), .IN2(n2590), .IN3(\regf[25][21] ), .IN4(n2410), 
        .Q(n868) );
  AO22X1 U894 ( .IN1(n2414), .IN2(n2593), .IN3(\regf[25][22] ), .IN4(n2410), 
        .Q(n869) );
  AO22X1 U895 ( .IN1(n2413), .IN2(n2596), .IN3(\regf[25][23] ), .IN4(n2410), 
        .Q(n870) );
  AO22X1 U896 ( .IN1(n2414), .IN2(n2599), .IN3(\regf[25][24] ), .IN4(n2410), 
        .Q(n871) );
  AO22X1 U897 ( .IN1(n2414), .IN2(n2602), .IN3(\regf[25][25] ), .IN4(n2410), 
        .Q(n872) );
  AO22X1 U898 ( .IN1(n2414), .IN2(n2605), .IN3(\regf[25][26] ), .IN4(n2410), 
        .Q(n873) );
  AO22X1 U899 ( .IN1(n2414), .IN2(n2608), .IN3(\regf[25][27] ), .IN4(n2410), 
        .Q(n874) );
  AO22X1 U900 ( .IN1(n2414), .IN2(n2611), .IN3(\regf[25][28] ), .IN4(n2410), 
        .Q(n875) );
  AO22X1 U901 ( .IN1(n2414), .IN2(n2614), .IN3(\regf[25][29] ), .IN4(n2410), 
        .Q(n876) );
  AO22X1 U902 ( .IN1(n2414), .IN2(n2617), .IN3(\regf[25][30] ), .IN4(n2410), 
        .Q(n877) );
  AO22X1 U903 ( .IN1(n2414), .IN2(n2620), .IN3(\regf[25][31] ), .IN4(n2410), 
        .Q(n878) );
  NOR3X0 U904 ( .IN1(wr_addr[1]), .IN2(wr_addr[2]), .IN3(n2714), .QN(n38) );
  AO22X1 U905 ( .IN1(n2407), .IN2(n2527), .IN3(\regf[26][0] ), .IN4(n2406), 
        .Q(n879) );
  AO22X1 U906 ( .IN1(n2407), .IN2(n2530), .IN3(\regf[26][1] ), .IN4(n2406), 
        .Q(n880) );
  AO22X1 U907 ( .IN1(n2407), .IN2(n2533), .IN3(\regf[26][2] ), .IN4(n2406), 
        .Q(n881) );
  AO22X1 U908 ( .IN1(n2407), .IN2(n2536), .IN3(\regf[26][3] ), .IN4(n2406), 
        .Q(n882) );
  AO22X1 U909 ( .IN1(n2408), .IN2(n2539), .IN3(\regf[26][4] ), .IN4(n2406), 
        .Q(n883) );
  AO22X1 U910 ( .IN1(n2409), .IN2(n2542), .IN3(\regf[26][5] ), .IN4(n2406), 
        .Q(n884) );
  AO22X1 U911 ( .IN1(n2408), .IN2(n2545), .IN3(\regf[26][6] ), .IN4(n2406), 
        .Q(n885) );
  AO22X1 U912 ( .IN1(n2408), .IN2(n2548), .IN3(\regf[26][7] ), .IN4(n2406), 
        .Q(n886) );
  AO22X1 U913 ( .IN1(n2409), .IN2(n2551), .IN3(\regf[26][8] ), .IN4(n2406), 
        .Q(n887) );
  AO22X1 U914 ( .IN1(n2409), .IN2(n2554), .IN3(\regf[26][9] ), .IN4(n2406), 
        .Q(n888) );
  AO22X1 U915 ( .IN1(n2408), .IN2(n2557), .IN3(\regf[26][10] ), .IN4(n2406), 
        .Q(n889) );
  AO22X1 U916 ( .IN1(n2408), .IN2(n2560), .IN3(\regf[26][11] ), .IN4(n2406), 
        .Q(n890) );
  AO22X1 U917 ( .IN1(n2408), .IN2(n2563), .IN3(\regf[26][12] ), .IN4(n2406), 
        .Q(n891) );
  AO22X1 U918 ( .IN1(n2408), .IN2(n2566), .IN3(\regf[26][13] ), .IN4(n2405), 
        .Q(n892) );
  AO22X1 U919 ( .IN1(n2408), .IN2(n2569), .IN3(\regf[26][14] ), .IN4(n73), .Q(
        n893) );
  AO22X1 U920 ( .IN1(n2408), .IN2(n2572), .IN3(\regf[26][15] ), .IN4(n73), .Q(
        n894) );
  AO22X1 U921 ( .IN1(n2408), .IN2(n2575), .IN3(\regf[26][16] ), .IN4(n73), .Q(
        n895) );
  AO22X1 U922 ( .IN1(n2408), .IN2(n2578), .IN3(\regf[26][17] ), .IN4(n73), .Q(
        n896) );
  AO22X1 U923 ( .IN1(n2409), .IN2(n2581), .IN3(\regf[26][18] ), .IN4(n73), .Q(
        n897) );
  AO22X1 U924 ( .IN1(n2408), .IN2(n2584), .IN3(\regf[26][19] ), .IN4(n73), .Q(
        n898) );
  AO22X1 U925 ( .IN1(n2409), .IN2(n2587), .IN3(\regf[26][20] ), .IN4(n2405), 
        .Q(n899) );
  AO22X1 U926 ( .IN1(n2408), .IN2(n2590), .IN3(\regf[26][21] ), .IN4(n2405), 
        .Q(n900) );
  AO22X1 U927 ( .IN1(n2409), .IN2(n2593), .IN3(\regf[26][22] ), .IN4(n2405), 
        .Q(n901) );
  AO22X1 U928 ( .IN1(n2408), .IN2(n2596), .IN3(\regf[26][23] ), .IN4(n2405), 
        .Q(n902) );
  AO22X1 U929 ( .IN1(n2409), .IN2(n2599), .IN3(\regf[26][24] ), .IN4(n2405), 
        .Q(n903) );
  AO22X1 U930 ( .IN1(n2409), .IN2(n2602), .IN3(\regf[26][25] ), .IN4(n2405), 
        .Q(n904) );
  AO22X1 U931 ( .IN1(n2409), .IN2(n2605), .IN3(\regf[26][26] ), .IN4(n2405), 
        .Q(n905) );
  AO22X1 U932 ( .IN1(n2409), .IN2(n2608), .IN3(\regf[26][27] ), .IN4(n2405), 
        .Q(n906) );
  AO22X1 U933 ( .IN1(n2409), .IN2(n2611), .IN3(\regf[26][28] ), .IN4(n2405), 
        .Q(n907) );
  AO22X1 U934 ( .IN1(n2409), .IN2(n2614), .IN3(\regf[26][29] ), .IN4(n2405), 
        .Q(n908) );
  AO22X1 U935 ( .IN1(n2409), .IN2(n2617), .IN3(\regf[26][30] ), .IN4(n2405), 
        .Q(n909) );
  AO22X1 U936 ( .IN1(n2409), .IN2(n2620), .IN3(\regf[26][31] ), .IN4(n2405), 
        .Q(n910) );
  NOR3X0 U937 ( .IN1(wr_addr[0]), .IN2(wr_addr[2]), .IN3(n2713), .QN(n41) );
  AO22X1 U938 ( .IN1(n2402), .IN2(n2527), .IN3(\regf[27][0] ), .IN4(n2401), 
        .Q(n911) );
  AO22X1 U939 ( .IN1(n2402), .IN2(n2530), .IN3(\regf[27][1] ), .IN4(n2401), 
        .Q(n912) );
  AO22X1 U940 ( .IN1(n2402), .IN2(n2533), .IN3(\regf[27][2] ), .IN4(n2401), 
        .Q(n913) );
  AO22X1 U941 ( .IN1(n2402), .IN2(n2536), .IN3(\regf[27][3] ), .IN4(n2401), 
        .Q(n914) );
  AO22X1 U942 ( .IN1(n2404), .IN2(n2539), .IN3(\regf[27][4] ), .IN4(n2401), 
        .Q(n915) );
  AO22X1 U943 ( .IN1(n2403), .IN2(n2542), .IN3(\regf[27][5] ), .IN4(n2401), 
        .Q(n916) );
  AO22X1 U944 ( .IN1(n2403), .IN2(n2545), .IN3(\regf[27][6] ), .IN4(n2401), 
        .Q(n917) );
  AO22X1 U945 ( .IN1(n2404), .IN2(n2548), .IN3(\regf[27][7] ), .IN4(n2401), 
        .Q(n918) );
  AO22X1 U946 ( .IN1(n2403), .IN2(n2551), .IN3(\regf[27][8] ), .IN4(n2401), 
        .Q(n919) );
  AO22X1 U947 ( .IN1(n2403), .IN2(n2554), .IN3(\regf[27][9] ), .IN4(n2401), 
        .Q(n920) );
  AO22X1 U948 ( .IN1(n2404), .IN2(n2557), .IN3(\regf[27][10] ), .IN4(n2401), 
        .Q(n921) );
  AO22X1 U949 ( .IN1(n2404), .IN2(n2560), .IN3(\regf[27][11] ), .IN4(n2401), 
        .Q(n922) );
  AO22X1 U950 ( .IN1(n2403), .IN2(n2563), .IN3(\regf[27][12] ), .IN4(n2401), 
        .Q(n923) );
  AO22X1 U951 ( .IN1(n2404), .IN2(n2566), .IN3(\regf[27][13] ), .IN4(n2400), 
        .Q(n924) );
  AO22X1 U952 ( .IN1(n2403), .IN2(n2569), .IN3(\regf[27][14] ), .IN4(n74), .Q(
        n925) );
  AO22X1 U953 ( .IN1(n2404), .IN2(n2572), .IN3(\regf[27][15] ), .IN4(n74), .Q(
        n926) );
  AO22X1 U954 ( .IN1(n2403), .IN2(n2575), .IN3(\regf[27][16] ), .IN4(n74), .Q(
        n927) );
  AO22X1 U955 ( .IN1(n2404), .IN2(n2578), .IN3(\regf[27][17] ), .IN4(n74), .Q(
        n928) );
  AO22X1 U956 ( .IN1(n2403), .IN2(n2581), .IN3(\regf[27][18] ), .IN4(n74), .Q(
        n929) );
  AO22X1 U957 ( .IN1(n2403), .IN2(n2584), .IN3(\regf[27][19] ), .IN4(n74), .Q(
        n930) );
  AO22X1 U958 ( .IN1(n2403), .IN2(n2587), .IN3(\regf[27][20] ), .IN4(n2400), 
        .Q(n931) );
  AO22X1 U959 ( .IN1(n2403), .IN2(n2590), .IN3(\regf[27][21] ), .IN4(n2400), 
        .Q(n932) );
  AO22X1 U960 ( .IN1(n2403), .IN2(n2593), .IN3(\regf[27][22] ), .IN4(n2400), 
        .Q(n933) );
  AO22X1 U961 ( .IN1(n2403), .IN2(n2596), .IN3(\regf[27][23] ), .IN4(n2400), 
        .Q(n934) );
  AO22X1 U962 ( .IN1(n2403), .IN2(n2599), .IN3(\regf[27][24] ), .IN4(n2400), 
        .Q(n935) );
  AO22X1 U963 ( .IN1(n2404), .IN2(n2602), .IN3(\regf[27][25] ), .IN4(n2400), 
        .Q(n936) );
  AO22X1 U964 ( .IN1(n2404), .IN2(n2605), .IN3(\regf[27][26] ), .IN4(n2400), 
        .Q(n937) );
  AO22X1 U965 ( .IN1(n2404), .IN2(n2608), .IN3(\regf[27][27] ), .IN4(n2400), 
        .Q(n938) );
  AO22X1 U966 ( .IN1(n2404), .IN2(n2611), .IN3(\regf[27][28] ), .IN4(n2400), 
        .Q(n939) );
  AO22X1 U967 ( .IN1(n2404), .IN2(n2614), .IN3(\regf[27][29] ), .IN4(n2400), 
        .Q(n940) );
  AO22X1 U968 ( .IN1(n2404), .IN2(n2617), .IN3(\regf[27][30] ), .IN4(n2400), 
        .Q(n941) );
  AO22X1 U969 ( .IN1(n2404), .IN2(n2620), .IN3(\regf[27][31] ), .IN4(n2400), 
        .Q(n942) );
  NOR3X0 U970 ( .IN1(n2714), .IN2(wr_addr[2]), .IN3(n2713), .QN(n43) );
  AO22X1 U971 ( .IN1(n2399), .IN2(n2527), .IN3(\regf[28][0] ), .IN4(n2397), 
        .Q(n943) );
  AO22X1 U972 ( .IN1(n2398), .IN2(n2530), .IN3(\regf[28][1] ), .IN4(n2397), 
        .Q(n944) );
  AO22X1 U973 ( .IN1(n2399), .IN2(n2533), .IN3(\regf[28][2] ), .IN4(n2397), 
        .Q(n945) );
  AO22X1 U974 ( .IN1(n2398), .IN2(n2536), .IN3(\regf[28][3] ), .IN4(n2397), 
        .Q(n946) );
  AO22X1 U975 ( .IN1(n2398), .IN2(n2539), .IN3(\regf[28][4] ), .IN4(n2397), 
        .Q(n947) );
  AO22X1 U976 ( .IN1(n2399), .IN2(n2542), .IN3(\regf[28][5] ), .IN4(n2397), 
        .Q(n948) );
  AO22X1 U977 ( .IN1(n2398), .IN2(n2545), .IN3(\regf[28][6] ), .IN4(n2397), 
        .Q(n949) );
  AO22X1 U978 ( .IN1(n2398), .IN2(n2548), .IN3(\regf[28][7] ), .IN4(n2397), 
        .Q(n950) );
  AO22X1 U979 ( .IN1(n2399), .IN2(n2551), .IN3(\regf[28][8] ), .IN4(n2397), 
        .Q(n951) );
  AO22X1 U980 ( .IN1(n2399), .IN2(n2554), .IN3(\regf[28][9] ), .IN4(n2397), 
        .Q(n952) );
  AO22X1 U981 ( .IN1(n2398), .IN2(n2557), .IN3(\regf[28][10] ), .IN4(n2397), 
        .Q(n953) );
  AO22X1 U982 ( .IN1(n2398), .IN2(n2560), .IN3(\regf[28][11] ), .IN4(n2397), 
        .Q(n954) );
  AO22X1 U983 ( .IN1(n2398), .IN2(n2563), .IN3(\regf[28][12] ), .IN4(n2397), 
        .Q(n955) );
  AO22X1 U984 ( .IN1(n2398), .IN2(n2566), .IN3(\regf[28][13] ), .IN4(n2396), 
        .Q(n956) );
  AO22X1 U985 ( .IN1(n2398), .IN2(n2569), .IN3(\regf[28][14] ), .IN4(n75), .Q(
        n957) );
  AO22X1 U986 ( .IN1(n2398), .IN2(n2572), .IN3(\regf[28][15] ), .IN4(n75), .Q(
        n958) );
  AO22X1 U987 ( .IN1(n2398), .IN2(n2575), .IN3(\regf[28][16] ), .IN4(n75), .Q(
        n959) );
  AO22X1 U988 ( .IN1(n2398), .IN2(n2578), .IN3(\regf[28][17] ), .IN4(n75), .Q(
        n960) );
  AO22X1 U989 ( .IN1(n2399), .IN2(n2581), .IN3(\regf[28][18] ), .IN4(n75), .Q(
        n961) );
  AO22X1 U990 ( .IN1(n2398), .IN2(n2584), .IN3(\regf[28][19] ), .IN4(n75), .Q(
        n962) );
  AO22X1 U991 ( .IN1(n2399), .IN2(n2587), .IN3(\regf[28][20] ), .IN4(n2396), 
        .Q(n963) );
  AO22X1 U992 ( .IN1(n2398), .IN2(n2590), .IN3(\regf[28][21] ), .IN4(n2396), 
        .Q(n964) );
  AO22X1 U993 ( .IN1(n2399), .IN2(n2593), .IN3(\regf[28][22] ), .IN4(n2396), 
        .Q(n965) );
  AO22X1 U994 ( .IN1(n2398), .IN2(n2596), .IN3(\regf[28][23] ), .IN4(n2396), 
        .Q(n966) );
  AO22X1 U995 ( .IN1(n2399), .IN2(n2599), .IN3(\regf[28][24] ), .IN4(n2396), 
        .Q(n967) );
  AO22X1 U996 ( .IN1(n2399), .IN2(n2602), .IN3(\regf[28][25] ), .IN4(n2396), 
        .Q(n968) );
  AO22X1 U997 ( .IN1(n2399), .IN2(n2605), .IN3(\regf[28][26] ), .IN4(n2396), 
        .Q(n969) );
  AO22X1 U998 ( .IN1(n2399), .IN2(n2608), .IN3(\regf[28][27] ), .IN4(n2396), 
        .Q(n970) );
  AO22X1 U999 ( .IN1(n2399), .IN2(n2611), .IN3(\regf[28][28] ), .IN4(n2396), 
        .Q(n971) );
  AO22X1 U1000 ( .IN1(n2399), .IN2(n2614), .IN3(\regf[28][29] ), .IN4(n2396), 
        .Q(n972) );
  AO22X1 U1001 ( .IN1(n2399), .IN2(n2617), .IN3(\regf[28][30] ), .IN4(n2396), 
        .Q(n973) );
  AO22X1 U1002 ( .IN1(n2399), .IN2(n2620), .IN3(\regf[28][31] ), .IN4(n2396), 
        .Q(n974) );
  AND3X1 U1003 ( .IN1(n2714), .IN2(n2713), .IN3(wr_addr[2]), .Q(n45) );
  AO22X1 U1004 ( .IN1(n2395), .IN2(n2527), .IN3(\regf[29][0] ), .IN4(n2393), 
        .Q(n975) );
  AO22X1 U1005 ( .IN1(n2394), .IN2(n2530), .IN3(\regf[29][1] ), .IN4(n2393), 
        .Q(n976) );
  AO22X1 U1006 ( .IN1(n2395), .IN2(n2533), .IN3(\regf[29][2] ), .IN4(n2393), 
        .Q(n977) );
  AO22X1 U1007 ( .IN1(n2394), .IN2(n2536), .IN3(\regf[29][3] ), .IN4(n2393), 
        .Q(n978) );
  AO22X1 U1008 ( .IN1(n2394), .IN2(n2539), .IN3(\regf[29][4] ), .IN4(n2393), 
        .Q(n979) );
  AO22X1 U1009 ( .IN1(n2395), .IN2(n2542), .IN3(\regf[29][5] ), .IN4(n2393), 
        .Q(n980) );
  AO22X1 U1010 ( .IN1(n2394), .IN2(n2545), .IN3(\regf[29][6] ), .IN4(n2393), 
        .Q(n981) );
  AO22X1 U1011 ( .IN1(n2394), .IN2(n2548), .IN3(\regf[29][7] ), .IN4(n2393), 
        .Q(n982) );
  AO22X1 U1012 ( .IN1(n2395), .IN2(n2551), .IN3(\regf[29][8] ), .IN4(n2393), 
        .Q(n983) );
  AO22X1 U1013 ( .IN1(n2395), .IN2(n2554), .IN3(\regf[29][9] ), .IN4(n2393), 
        .Q(n984) );
  AO22X1 U1014 ( .IN1(n2394), .IN2(n2557), .IN3(\regf[29][10] ), .IN4(n2393), 
        .Q(n985) );
  AO22X1 U1015 ( .IN1(n2394), .IN2(n2560), .IN3(\regf[29][11] ), .IN4(n2393), 
        .Q(n986) );
  AO22X1 U1016 ( .IN1(n2394), .IN2(n2563), .IN3(\regf[29][12] ), .IN4(n2393), 
        .Q(n987) );
  AO22X1 U1017 ( .IN1(n2394), .IN2(n2566), .IN3(\regf[29][13] ), .IN4(n2392), 
        .Q(n988) );
  AO22X1 U1018 ( .IN1(n2394), .IN2(n2569), .IN3(\regf[29][14] ), .IN4(n76), 
        .Q(n989) );
  AO22X1 U1019 ( .IN1(n2394), .IN2(n2572), .IN3(\regf[29][15] ), .IN4(n76), 
        .Q(n990) );
  AO22X1 U1020 ( .IN1(n2394), .IN2(n2575), .IN3(\regf[29][16] ), .IN4(n76), 
        .Q(n991) );
  AO22X1 U1021 ( .IN1(n2394), .IN2(n2578), .IN3(\regf[29][17] ), .IN4(n76), 
        .Q(n992) );
  AO22X1 U1022 ( .IN1(n2395), .IN2(n2581), .IN3(\regf[29][18] ), .IN4(n76), 
        .Q(n993) );
  AO22X1 U1023 ( .IN1(n2394), .IN2(n2584), .IN3(\regf[29][19] ), .IN4(n76), 
        .Q(n994) );
  AO22X1 U1024 ( .IN1(n2395), .IN2(n2587), .IN3(\regf[29][20] ), .IN4(n2392), 
        .Q(n995) );
  AO22X1 U1025 ( .IN1(n2394), .IN2(n2590), .IN3(\regf[29][21] ), .IN4(n2392), 
        .Q(n996) );
  AO22X1 U1026 ( .IN1(n2395), .IN2(n2593), .IN3(\regf[29][22] ), .IN4(n2392), 
        .Q(n997) );
  AO22X1 U1027 ( .IN1(n2394), .IN2(n2596), .IN3(\regf[29][23] ), .IN4(n2392), 
        .Q(n998) );
  AO22X1 U1028 ( .IN1(n2395), .IN2(n2599), .IN3(\regf[29][24] ), .IN4(n2392), 
        .Q(n999) );
  AO22X1 U1029 ( .IN1(n2395), .IN2(n2602), .IN3(\regf[29][25] ), .IN4(n2392), 
        .Q(n1000) );
  AO22X1 U1030 ( .IN1(n2395), .IN2(n2605), .IN3(\regf[29][26] ), .IN4(n2392), 
        .Q(n1001) );
  AO22X1 U1031 ( .IN1(n2395), .IN2(n2608), .IN3(\regf[29][27] ), .IN4(n2392), 
        .Q(n1002) );
  AO22X1 U1032 ( .IN1(n2395), .IN2(n2611), .IN3(\regf[29][28] ), .IN4(n2392), 
        .Q(n1003) );
  AO22X1 U1033 ( .IN1(n2395), .IN2(n2614), .IN3(\regf[29][29] ), .IN4(n2392), 
        .Q(n1004) );
  AO22X1 U1034 ( .IN1(n2395), .IN2(n2617), .IN3(\regf[29][30] ), .IN4(n2392), 
        .Q(n1005) );
  AO22X1 U1035 ( .IN1(n2395), .IN2(n2620), .IN3(\regf[29][31] ), .IN4(n2392), 
        .Q(n1006) );
  AND3X1 U1036 ( .IN1(wr_addr[0]), .IN2(n2713), .IN3(wr_addr[2]), .Q(n47) );
  AO22X1 U1037 ( .IN1(n2391), .IN2(n2527), .IN3(\regf[30][0] ), .IN4(n2389), 
        .Q(n1007) );
  AO22X1 U1038 ( .IN1(n2390), .IN2(n2530), .IN3(\regf[30][1] ), .IN4(n2389), 
        .Q(n1008) );
  AO22X1 U1039 ( .IN1(n2391), .IN2(n2533), .IN3(\regf[30][2] ), .IN4(n2389), 
        .Q(n1009) );
  AO22X1 U1040 ( .IN1(n2390), .IN2(n2536), .IN3(\regf[30][3] ), .IN4(n2389), 
        .Q(n1010) );
  AO22X1 U1041 ( .IN1(n2390), .IN2(n2539), .IN3(\regf[30][4] ), .IN4(n2389), 
        .Q(n1011) );
  AO22X1 U1042 ( .IN1(n2391), .IN2(n2542), .IN3(\regf[30][5] ), .IN4(n2389), 
        .Q(n1012) );
  AO22X1 U1043 ( .IN1(n2390), .IN2(n2545), .IN3(\regf[30][6] ), .IN4(n2389), 
        .Q(n1013) );
  AO22X1 U1044 ( .IN1(n2390), .IN2(n2548), .IN3(\regf[30][7] ), .IN4(n2389), 
        .Q(n1014) );
  AO22X1 U1045 ( .IN1(n2391), .IN2(n2551), .IN3(\regf[30][8] ), .IN4(n2389), 
        .Q(n1015) );
  AO22X1 U1046 ( .IN1(n2391), .IN2(n2554), .IN3(\regf[30][9] ), .IN4(n2389), 
        .Q(n1016) );
  AO22X1 U1047 ( .IN1(n2390), .IN2(n2557), .IN3(\regf[30][10] ), .IN4(n2389), 
        .Q(n1017) );
  AO22X1 U1048 ( .IN1(n2390), .IN2(n2560), .IN3(\regf[30][11] ), .IN4(n2389), 
        .Q(n1018) );
  AO22X1 U1049 ( .IN1(n2390), .IN2(n2563), .IN3(\regf[30][12] ), .IN4(n2389), 
        .Q(n1019) );
  AO22X1 U1050 ( .IN1(n2390), .IN2(n2566), .IN3(\regf[30][13] ), .IN4(n2388), 
        .Q(n1020) );
  AO22X1 U1051 ( .IN1(n2390), .IN2(n2569), .IN3(\regf[30][14] ), .IN4(n77), 
        .Q(n1021) );
  AO22X1 U1052 ( .IN1(n2390), .IN2(n2572), .IN3(\regf[30][15] ), .IN4(n77), 
        .Q(n1022) );
  AO22X1 U1053 ( .IN1(n2390), .IN2(n2575), .IN3(\regf[30][16] ), .IN4(n77), 
        .Q(n1023) );
  AO22X1 U1054 ( .IN1(n2390), .IN2(n2578), .IN3(\regf[30][17] ), .IN4(n77), 
        .Q(n1024) );
  AO22X1 U1055 ( .IN1(n2391), .IN2(n2581), .IN3(\regf[30][18] ), .IN4(n77), 
        .Q(n1025) );
  AO22X1 U1056 ( .IN1(n2390), .IN2(n2584), .IN3(\regf[30][19] ), .IN4(n77), 
        .Q(n1026) );
  AO22X1 U1057 ( .IN1(n2391), .IN2(n2587), .IN3(\regf[30][20] ), .IN4(n2388), 
        .Q(n1027) );
  AO22X1 U1058 ( .IN1(n2390), .IN2(n2590), .IN3(\regf[30][21] ), .IN4(n2388), 
        .Q(n1028) );
  AO22X1 U1059 ( .IN1(n2391), .IN2(n2593), .IN3(\regf[30][22] ), .IN4(n2388), 
        .Q(n1029) );
  AO22X1 U1060 ( .IN1(n2390), .IN2(n2596), .IN3(\regf[30][23] ), .IN4(n2388), 
        .Q(n1030) );
  AO22X1 U1061 ( .IN1(n2391), .IN2(n2599), .IN3(\regf[30][24] ), .IN4(n2388), 
        .Q(n1031) );
  AO22X1 U1062 ( .IN1(n2391), .IN2(n2602), .IN3(\regf[30][25] ), .IN4(n2388), 
        .Q(n1032) );
  AO22X1 U1063 ( .IN1(n2391), .IN2(n2605), .IN3(\regf[30][26] ), .IN4(n2388), 
        .Q(n1033) );
  AO22X1 U1064 ( .IN1(n2391), .IN2(n2608), .IN3(\regf[30][27] ), .IN4(n2388), 
        .Q(n1034) );
  AO22X1 U1065 ( .IN1(n2391), .IN2(n2611), .IN3(\regf[30][28] ), .IN4(n2388), 
        .Q(n1035) );
  AO22X1 U1066 ( .IN1(n2391), .IN2(n2614), .IN3(\regf[30][29] ), .IN4(n2388), 
        .Q(n1036) );
  AO22X1 U1067 ( .IN1(n2391), .IN2(n2617), .IN3(\regf[30][30] ), .IN4(n2388), 
        .Q(n1037) );
  AO22X1 U1068 ( .IN1(n2391), .IN2(n2620), .IN3(\regf[30][31] ), .IN4(n2388), 
        .Q(n1038) );
  AND3X1 U1069 ( .IN1(wr_addr[1]), .IN2(n2714), .IN3(wr_addr[2]), .Q(n49) );
  AO22X1 U1070 ( .IN1(n2387), .IN2(n2527), .IN3(\regf[31][0] ), .IN4(n2385), 
        .Q(n1039) );
  AO22X1 U1071 ( .IN1(n2386), .IN2(n2530), .IN3(\regf[31][1] ), .IN4(n2385), 
        .Q(n1040) );
  AO22X1 U1072 ( .IN1(n2387), .IN2(n2533), .IN3(\regf[31][2] ), .IN4(n2385), 
        .Q(n1041) );
  AO22X1 U1073 ( .IN1(n2386), .IN2(n2536), .IN3(\regf[31][3] ), .IN4(n2385), 
        .Q(n1042) );
  AO22X1 U1074 ( .IN1(n2386), .IN2(n2539), .IN3(\regf[31][4] ), .IN4(n2385), 
        .Q(n1043) );
  AO22X1 U1075 ( .IN1(n2387), .IN2(n2542), .IN3(\regf[31][5] ), .IN4(n2385), 
        .Q(n1044) );
  AO22X1 U1076 ( .IN1(n2386), .IN2(n2545), .IN3(\regf[31][6] ), .IN4(n2385), 
        .Q(n1045) );
  AO22X1 U1077 ( .IN1(n2386), .IN2(n2548), .IN3(\regf[31][7] ), .IN4(n2385), 
        .Q(n1046) );
  AO22X1 U1078 ( .IN1(n2387), .IN2(n2551), .IN3(\regf[31][8] ), .IN4(n2385), 
        .Q(n1047) );
  AO22X1 U1079 ( .IN1(n2387), .IN2(n2554), .IN3(\regf[31][9] ), .IN4(n2385), 
        .Q(n1048) );
  AO22X1 U1080 ( .IN1(n2386), .IN2(n2557), .IN3(\regf[31][10] ), .IN4(n2385), 
        .Q(n1049) );
  AO22X1 U1081 ( .IN1(n2386), .IN2(n2560), .IN3(\regf[31][11] ), .IN4(n2385), 
        .Q(n1050) );
  AO22X1 U1082 ( .IN1(n2386), .IN2(n2563), .IN3(\regf[31][12] ), .IN4(n2385), 
        .Q(n1051) );
  AO22X1 U1083 ( .IN1(n2386), .IN2(n2566), .IN3(\regf[31][13] ), .IN4(n2384), 
        .Q(n1052) );
  AO22X1 U1084 ( .IN1(n2386), .IN2(n2569), .IN3(\regf[31][14] ), .IN4(n78), 
        .Q(n1053) );
  AO22X1 U1085 ( .IN1(n2386), .IN2(n2572), .IN3(\regf[31][15] ), .IN4(n78), 
        .Q(n1054) );
  AO22X1 U1086 ( .IN1(n2386), .IN2(n2575), .IN3(\regf[31][16] ), .IN4(n78), 
        .Q(n1055) );
  AO22X1 U1087 ( .IN1(n2386), .IN2(n2578), .IN3(\regf[31][17] ), .IN4(n78), 
        .Q(n1056) );
  AO22X1 U1088 ( .IN1(n2387), .IN2(n2581), .IN3(\regf[31][18] ), .IN4(n78), 
        .Q(n1057) );
  AO22X1 U1089 ( .IN1(n2386), .IN2(n2584), .IN3(\regf[31][19] ), .IN4(n78), 
        .Q(n1058) );
  AO22X1 U1090 ( .IN1(n2387), .IN2(n2587), .IN3(\regf[31][20] ), .IN4(n2384), 
        .Q(n1059) );
  AO22X1 U1091 ( .IN1(n2386), .IN2(n2590), .IN3(\regf[31][21] ), .IN4(n2384), 
        .Q(n1060) );
  AO22X1 U1092 ( .IN1(n2387), .IN2(n2593), .IN3(\regf[31][22] ), .IN4(n2384), 
        .Q(n1061) );
  AO22X1 U1093 ( .IN1(n2386), .IN2(n2596), .IN3(\regf[31][23] ), .IN4(n2384), 
        .Q(n1062) );
  AO22X1 U1094 ( .IN1(n2387), .IN2(n2599), .IN3(\regf[31][24] ), .IN4(n2384), 
        .Q(n1063) );
  AO22X1 U1095 ( .IN1(n2387), .IN2(n2602), .IN3(\regf[31][25] ), .IN4(n2384), 
        .Q(n1064) );
  AO22X1 U1096 ( .IN1(n2387), .IN2(n2605), .IN3(\regf[31][26] ), .IN4(n2384), 
        .Q(n1065) );
  AO22X1 U1097 ( .IN1(n2387), .IN2(n2608), .IN3(\regf[31][27] ), .IN4(n2384), 
        .Q(n1066) );
  AO22X1 U1098 ( .IN1(n2387), .IN2(n2611), .IN3(\regf[31][28] ), .IN4(n2384), 
        .Q(n1067) );
  AO22X1 U1099 ( .IN1(n2387), .IN2(n2614), .IN3(\regf[31][29] ), .IN4(n2384), 
        .Q(n1068) );
  AO22X1 U1100 ( .IN1(n2387), .IN2(n2617), .IN3(\regf[31][30] ), .IN4(n2384), 
        .Q(n1069) );
  AO22X1 U1101 ( .IN1(n2387), .IN2(n2620), .IN3(\regf[31][31] ), .IN4(n2384), 
        .Q(n1070) );
  AND3X1 U1102 ( .IN1(wr_addr[1]), .IN2(wr_addr[0]), .IN3(wr_addr[2]), .Q(n51)
         );
  AND3X1 U1103 ( .IN1(wr_addr[3]), .IN2(wr_en), .IN3(wr_addr[4]), .Q(n71) );
  NAND3X1 U1104 ( .IN1(\regf[3][31] ), .IN2(n1213), .IN3(n1376), .QN(n2233) );
  MUX21X1 U1105 ( .IN1(n1693), .IN2(n1688), .S(n1910), .Q(rd_dataA[24]) );
  MUX21X1 U1106 ( .IN1(n1713), .IN2(n1708), .S(n1910), .Q(rd_dataA[26]) );
  MUX41X2 U1107 ( .IN1(n2189), .IN3(n2187), .IN2(n2188), .IN4(n2186), .S0(
        n2379), .S1(n2373), .Q(n2190) );
  MUX41X2 U1108 ( .IN1(n1949), .IN3(n1947), .IN2(n1948), .IN4(n1946), .S0(
        n2375), .S1(n2369), .Q(n1950) );
  MUX21X2 U1109 ( .IN1(n1673), .IN2(n1668), .S(n1910), .Q(rd_dataA[22]) );
  MUX21X2 U1110 ( .IN1(n2050), .IN2(n2045), .S(n2381), .Q(rd_dataB[13]) );
  MUX21X2 U1111 ( .IN1(n2020), .IN2(n2015), .S(n2381), .Q(rd_dataB[10]) );
  MUX21X2 U1112 ( .IN1(n1553), .IN2(n1548), .S(n1909), .Q(rd_dataA[10]) );
  NAND3X1 U1113 ( .IN1(\regf[3][11] ), .IN2(n1297), .IN3(n1132), .QN(n1846) );
  MUX41X2 U1114 ( .IN1(n2179), .IN3(n2177), .IN2(n2178), .IN4(n2176), .S0(
        n2379), .S1(n2373), .Q(n2180) );
  MUX41X2 U1115 ( .IN1(n1722), .IN3(n1720), .IN2(n1721), .IN4(n1719), .S0(
        n1907), .S1(n1901), .Q(n1723) );
  MUX21X1 U1116 ( .IN1(n1950), .IN2(n1945), .S(n2380), .Q(rd_dataB[3]) );
  MUX21X2 U1117 ( .IN1(n1780), .IN2(n1781), .S(n1314), .Q(n1783) );
  MUX21X2 U1118 ( .IN1(n2230), .IN2(n2225), .S(n2382), .Q(rd_dataB[31]) );
  MUX21X2 U1119 ( .IN1(n2160), .IN2(n2155), .S(n2382), .Q(rd_dataB[24]) );
  MUX41X1 U1120 ( .IN1(n2159), .IN3(n2157), .IN2(n2158), .IN4(n2156), .S0(
        n2378), .S1(n2372), .Q(n2160) );
  INVX0 U1121 ( .INP(n2366), .ZN(n1071) );
  DELLN1X2 U1122 ( .INP(n1438), .Z(n1072) );
  DELLN1X2 U1123 ( .INP(n1400), .Z(n1073) );
  MUX21X2 U1124 ( .IN1(n1868), .IN2(n1869), .S(n1303), .Q(n1871) );
  MUX21X1 U1125 ( .IN1(n1503), .IN2(n1498), .S(n1908), .Q(rd_dataA[5]) );
  DELLN1X2 U1126 ( .INP(n1427), .Z(n1074) );
  NAND3X1 U1127 ( .IN1(\regf[3][31] ), .IN2(n1293), .IN3(n1427), .QN(n1766) );
  INVX0 U1128 ( .INP(n1413), .ZN(n1075) );
  INVX0 U1129 ( .INP(n1413), .ZN(n1076) );
  INVX0 U1130 ( .INP(n2366), .ZN(n1077) );
  INVX0 U1131 ( .INP(n2366), .ZN(n1078) );
  NAND3X1 U1132 ( .IN1(\regf[3][29] ), .IN2(n1215), .IN3(n1078), .QN(n2241) );
  DELLN1X2 U1133 ( .INP(n1398), .Z(n1079) );
  MUX41X2 U1134 ( .IN1(n1984), .IN3(n1982), .IN2(n1983), .IN4(n1981), .S0(
        n2375), .S1(n2369), .Q(n1985) );
  MUX41X2 U1135 ( .IN1(n2054), .IN3(n2052), .IN2(n2053), .IN4(n2051), .S0(
        n2377), .S1(n2371), .Q(n2055) );
  MUX41X2 U1136 ( .IN1(n2004), .IN3(n2002), .IN2(n2003), .IN4(n2001), .S0(
        n2376), .S1(n2370), .Q(n2005) );
  MUX21X1 U1137 ( .IN1(n1563), .IN2(n1558), .S(n1909), .Q(rd_dataA[11]) );
  MUX21X1 U1138 ( .IN1(n1513), .IN2(n1508), .S(n1908), .Q(rd_dataA[6]) );
  DELLN1X2 U1139 ( .INP(n1427), .Z(n1080) );
  NAND3X1 U1140 ( .IN1(\regf[3][6] ), .IN2(n1296), .IN3(n1398), .QN(n1866) );
  MUX41X2 U1141 ( .IN1(n2024), .IN3(n2022), .IN2(n2023), .IN4(n2021), .S0(
        n2376), .S1(n2370), .Q(n2025) );
  MUX21X2 U1142 ( .IN1(n1990), .IN2(n1985), .S(n2380), .Q(rd_dataB[7]) );
  MUX21X2 U1143 ( .IN1(n2060), .IN2(n2055), .S(n2381), .Q(rd_dataB[14]) );
  MUX21X2 U1144 ( .IN1(n2010), .IN2(n2005), .S(n2381), .Q(rd_dataB[9]) );
  MUX41X2 U1145 ( .IN1(n2124), .IN3(n2122), .IN2(n2123), .IN4(n2121), .S0(
        n2378), .S1(n2372), .Q(n2125) );
  MUX41X1 U1146 ( .IN1(n2069), .IN3(n2067), .IN2(n2068), .IN4(n2066), .S0(
        n2377), .S1(n2371), .Q(n2070) );
  MUX21X2 U1147 ( .IN1(n2210), .IN2(n2205), .S(n2382), .Q(rd_dataB[29]) );
  MUX21X2 U1148 ( .IN1(n1453), .IN2(n1448), .S(n1908), .Q(rd_dataA[0]) );
  MUX21X2 U1149 ( .IN1(n1613), .IN2(n1608), .S(n1909), .Q(rd_dataA[16]) );
  MUX21X2 U1150 ( .IN1(n1763), .IN2(n1758), .S(n1910), .Q(rd_dataA[31]) );
  MUX21X2 U1151 ( .IN1(n1703), .IN2(n1698), .S(n1910), .Q(rd_dataA[25]) );
  MUX41X2 U1152 ( .IN1(n1737), .IN3(n1735), .IN2(n1736), .IN4(n1734), .S0(
        n1907), .S1(n1901), .Q(n1738) );
  MUX41X2 U1153 ( .IN1(n1577), .IN3(n1575), .IN2(n1576), .IN4(n1574), .S0(
        n1904), .S1(n1898), .Q(n1578) );
  MUX41X2 U1154 ( .IN1(n1482), .IN3(n1480), .IN2(n1481), .IN4(n1479), .S0(
        n1903), .S1(n1897), .Q(n1483) );
  MUX41X1 U1155 ( .IN1(\regf[25][14] ), .IN3(\regf[27][14] ), .IN2(
        \regf[24][14] ), .IN4(\regf[26][14] ), .S0(n1334), .S1(n1083), .Q(
        n1585) );
  MUX21X2 U1156 ( .IN1(n1593), .IN2(n1588), .S(n1909), .Q(rd_dataA[14]) );
  MUX41X1 U1157 ( .IN1(n1587), .IN3(n1585), .IN2(n1586), .IN4(n1584), .S0(
        n1905), .S1(n1899), .Q(n1588) );
  DELLN1X2 U1158 ( .INP(n1442), .Z(n1081) );
  INVX0 U1159 ( .INP(n1893), .ZN(n1082) );
  INVX0 U1160 ( .INP(n1442), .ZN(n1083) );
  INVX0 U1161 ( .INP(n1415), .ZN(n1084) );
  INVX0 U1162 ( .INP(n1415), .ZN(n1085) );
  DELLN1X2 U1163 ( .INP(n1400), .Z(n1086) );
  INVX0 U1164 ( .INP(n1894), .ZN(n1087) );
  MUX21X1 U1165 ( .IN1(n2343), .IN2(n2344), .S(n1229), .Q(n2346) );
  NAND3X1 U1166 ( .IN1(\regf[3][8] ), .IN2(n1247), .IN3(n1386), .QN(n2325) );
  MUX41X1 U1167 ( .IN1(\regf[28][5] ), .IN3(\regf[30][5] ), .IN2(\regf[29][5] ), .IN4(\regf[31][5] ), .S0(n1328), .S1(n1419), .Q(n1494) );
  NAND3X1 U1168 ( .IN1(\regf[3][26] ), .IN2(n1302), .IN3(n1435), .QN(n1786) );
  MUX41X1 U1169 ( .IN1(\regf[4][26] ), .IN3(\regf[6][26] ), .IN2(\regf[5][26] ), .IN4(\regf[7][26] ), .S0(n1351), .S1(n1434), .Q(n1711) );
  MUX41X1 U1170 ( .IN1(\regf[28][29] ), .IN3(\regf[30][29] ), .IN2(
        \regf[29][29] ), .IN4(\regf[31][29] ), .S0(n1346), .S1(n1419), .Q(
        n1734) );
  MUX41X1 U1171 ( .IN1(\regf[20][30] ), .IN3(\regf[22][30] ), .IN2(
        \regf[21][30] ), .IN4(\regf[23][30] ), .S0(n1347), .S1(n1423), .Q(
        n1746) );
  MUX41X1 U1172 ( .IN1(\regf[16][31] ), .IN3(\regf[18][31] ), .IN2(
        \regf[17][31] ), .IN4(\regf[19][31] ), .S0(n1343), .S1(n1418), .Q(
        n1757) );
  MUX41X1 U1173 ( .IN1(n1969), .IN3(n1967), .IN2(n1968), .IN4(n1966), .S0(
        n2375), .S1(n2369), .Q(n1970) );
  MUX41X1 U1174 ( .IN1(n1979), .IN3(n1977), .IN2(n1978), .IN4(n1976), .S0(
        n2375), .S1(n2369), .Q(n1980) );
  MUX41X1 U1175 ( .IN1(n2049), .IN3(n2047), .IN2(n2048), .IN4(n2046), .S0(
        n2376), .S1(n2370), .Q(n2050) );
  MUX41X1 U1176 ( .IN1(n2084), .IN3(n2082), .IN2(n2083), .IN4(n2081), .S0(
        n2377), .S1(n2371), .Q(n2085) );
  MUX41X1 U1177 ( .IN1(\regf[20][11] ), .IN3(\regf[22][11] ), .IN2(
        \regf[21][11] ), .IN4(\regf[23][11] ), .S0(n1342), .S1(n1418), .Q(
        n1556) );
  NAND2X0 U1178 ( .IN1(n62), .IN2(n51), .QN(n69) );
  MUX21X2 U1179 ( .IN1(n1920), .IN2(n1915), .S(n2380), .Q(rd_dataB[0]) );
  MUX21X2 U1180 ( .IN1(n2110), .IN2(n2105), .S(n2381), .Q(rd_dataB[19]) );
  MUX41X2 U1181 ( .IN1(n2214), .IN3(n2212), .IN2(n2213), .IN4(n2211), .S0(
        n2379), .S1(n2373), .Q(n2215) );
  MUX21X2 U1182 ( .IN1(n2220), .IN2(n2215), .S(n2382), .Q(rd_dataB[30]) );
  MUX41X2 U1183 ( .IN1(n2029), .IN3(n2027), .IN2(n2028), .IN4(n2026), .S0(
        n2376), .S1(n2370), .Q(n2030) );
  MUX21X2 U1184 ( .IN1(n2311), .IN2(n2312), .S(n1232), .Q(n2314) );
  MUX41X1 U1185 ( .IN1(n2209), .IN3(n2207), .IN2(n2208), .IN4(n2206), .S0(
        n2379), .S1(n2373), .Q(n2210) );
  DELLN1X2 U1186 ( .INP(n1371), .Z(n1088) );
  DELLN1X2 U1187 ( .INP(n1371), .Z(n1089) );
  MUX21X2 U1188 ( .IN1(n2090), .IN2(n2085), .S(n2381), .Q(rd_dataB[17]) );
  INVX0 U1189 ( .INP(n2365), .ZN(n1090) );
  MUX21X2 U1190 ( .IN1(n2200), .IN2(n2195), .S(n2382), .Q(rd_dataB[28]) );
  DELLN1X2 U1191 ( .INP(n1400), .Z(n1091) );
  DELLN1X2 U1192 ( .INP(n1103), .Z(n1092) );
  MUX21X2 U1193 ( .IN1(n1940), .IN2(n1935), .S(n2380), .Q(rd_dataB[2]) );
  MUX21X2 U1194 ( .IN1(n1960), .IN2(n1955), .S(n2380), .Q(rd_dataB[4]) );
  DELLN1X2 U1195 ( .INP(n1380), .Z(n1093) );
  DELLN1X2 U1196 ( .INP(n1378), .Z(n1094) );
  DELLN1X2 U1197 ( .INP(n1378), .Z(n1095) );
  DELLN1X2 U1198 ( .INP(n1371), .Z(n1096) );
  NAND3X1 U1199 ( .IN1(\regf[3][16] ), .IN2(n1292), .IN3(n1400), .QN(n1826) );
  INVX0 U1200 ( .INP(n2366), .ZN(n1097) );
  MUX21X2 U1201 ( .IN1(n2100), .IN2(n2095), .S(n2381), .Q(rd_dataB[18]) );
  OR2X1 U1202 ( .IN1(n1098), .IN2(n1355), .Q(n2256) );
  MUX21X2 U1203 ( .IN1(n2170), .IN2(n2165), .S(n2382), .Q(rd_dataB[25]) );
  MUX41X1 U1204 ( .IN1(n2169), .IN3(n2167), .IN2(n2168), .IN4(n2166), .S0(
        n2378), .S1(n2372), .Q(n2170) );
  OR2X1 U1205 ( .IN1(n1099), .IN2(n1382), .Q(n2344) );
  MUX21X2 U1206 ( .IN1(n1733), .IN2(n1728), .S(n1910), .Q(rd_dataA[28]) );
  MUX21X2 U1207 ( .IN1(n1633), .IN2(n1628), .S(n1909), .Q(rd_dataA[18]) );
  MUX41X2 U1208 ( .IN1(n1994), .IN3(n1992), .IN2(n1993), .IN4(n1991), .S0(
        n2376), .S1(n2370), .Q(n1995) );
  MUX21X2 U1209 ( .IN1(n2255), .IN2(n2256), .S(n1216), .Q(n2258) );
  MUX21X2 U1210 ( .IN1(n2315), .IN2(n2316), .S(n1234), .Q(n2318) );
  MUX21X2 U1211 ( .IN1(n2331), .IN2(n2332), .S(n1227), .Q(n2334) );
  MUX21X2 U1212 ( .IN1(n1643), .IN2(n1638), .S(n1909), .Q(rd_dataA[19]) );
  MUX21X2 U1213 ( .IN1(n1753), .IN2(n1748), .S(n1910), .Q(rd_dataA[30]) );
  OR2X1 U1214 ( .IN1(n1100), .IN2(n1395), .Q(n2336) );
  MUX41X1 U1215 ( .IN1(\regf[20][18] ), .IN3(\regf[22][18] ), .IN2(
        \regf[21][18] ), .IN4(\regf[23][18] ), .S0(n1351), .S1(n1087), .Q(
        n1626) );
  INVX0 U1216 ( .INP(n1894), .ZN(n1101) );
  MUX21X2 U1217 ( .IN1(n2000), .IN2(n1995), .S(n2381), .Q(rd_dataB[8]) );
  OR2X1 U1218 ( .IN1(n1102), .IN2(n1397), .Q(n1885) );
  MUX41X1 U1219 ( .IN1(n1462), .IN3(n1460), .IN2(n1461), .IN4(n1459), .S0(
        n1902), .S1(n1896), .Q(n1463) );
  MUX21X2 U1220 ( .IN1(n1816), .IN2(n1817), .S(n1319), .Q(n1819) );
  MUX21X2 U1221 ( .IN1(n1812), .IN2(n1813), .S(n1309), .Q(n1815) );
  MUX21X2 U1222 ( .IN1(n1872), .IN2(n1873), .S(n1305), .Q(n1875) );
  MUX21X2 U1223 ( .IN1(n2335), .IN2(n2336), .S(n1224), .Q(n2338) );
  MUX41X2 U1224 ( .IN1(n1597), .IN3(n1595), .IN2(n1596), .IN4(n1594), .S0(
        n1905), .S1(n1899), .Q(n1598) );
  MUX41X1 U1225 ( .IN1(\regf[20][17] ), .IN3(\regf[22][17] ), .IN2(
        \regf[21][17] ), .IN4(\regf[23][17] ), .S0(n1345), .S1(n1409), .Q(
        n1616) );
  INVX0 U1226 ( .INP(n2360), .ZN(n1103) );
  MUX41X2 U1227 ( .IN1(n1537), .IN3(n1535), .IN2(n1536), .IN4(n1534), .S0(
        n1904), .S1(n1898), .Q(n1538) );
  MUX41X1 U1228 ( .IN1(\regf[16][26] ), .IN3(\regf[18][26] ), .IN2(
        \regf[17][26] ), .IN4(\regf[19][26] ), .S0(n1351), .S1(n1407), .Q(
        n1707) );
  NAND3X1 U1229 ( .IN1(\regf[3][29] ), .IN2(n1302), .IN3(n1407), .QN(n1774) );
  MUX21X2 U1230 ( .IN1(n1603), .IN2(n1598), .S(n1909), .Q(rd_dataA[15]) );
  MUX41X1 U1231 ( .IN1(\regf[12][19] ), .IN3(\regf[14][19] ), .IN2(
        \regf[13][19] ), .IN4(\regf[15][19] ), .S0(n1352), .S1(n1183), .Q(
        n1639) );
  MUX41X2 U1232 ( .IN1(n1617), .IN3(n1615), .IN2(n1616), .IN4(n1614), .S0(
        n1905), .S1(n1899), .Q(n1618) );
  MUX41X2 U1233 ( .IN1(n1657), .IN3(n1655), .IN2(n1656), .IN4(n1654), .S0(
        n1906), .S1(n1900), .Q(n1658) );
  DELLN1X2 U1234 ( .INP(n1388), .Z(n1104) );
  DELLN1X2 U1235 ( .INP(n1378), .Z(n1105) );
  INVX0 U1236 ( .INP(n2362), .ZN(n1106) );
  INVX0 U1237 ( .INP(n2361), .ZN(n1107) );
  DELLN1X2 U1238 ( .INP(n1427), .Z(n1108) );
  MUX41X1 U1239 ( .IN1(n1512), .IN3(n1510), .IN2(n1511), .IN4(n1509), .S0(
        n1903), .S1(n1897), .Q(n1513) );
  NAND3X2 U1240 ( .IN1(\regf[3][2] ), .IN2(n1205), .IN3(n1374), .QN(n2349) );
  MUX21X2 U1241 ( .IN1(n1623), .IN2(n1618), .S(n1909), .Q(rd_dataA[17]) );
  MUX21X2 U1242 ( .IN1(n1583), .IN2(n1578), .S(n1909), .Q(rd_dataA[13]) );
  MUX21X2 U1243 ( .IN1(n1663), .IN2(n1658), .S(n1910), .Q(rd_dataA[21]) );
  MUX21X2 U1244 ( .IN1(n1743), .IN2(n1738), .S(n1910), .Q(rd_dataA[29]) );
  MUX21X2 U1245 ( .IN1(n1573), .IN2(n1568), .S(n1909), .Q(rd_dataA[12]) );
  MUX41X1 U1246 ( .IN1(\regf[12][2] ), .IN3(\regf[14][2] ), .IN2(\regf[13][2] ), .IN4(\regf[15][2] ), .S0(n1351), .S1(n1108), .Q(n1469) );
  MUX41X1 U1247 ( .IN1(\regf[20][0] ), .IN3(\regf[22][0] ), .IN2(\regf[21][0] ), .IN4(\regf[23][0] ), .S0(n1348), .S1(n1108), .Q(n1446) );
  INVX0 U1248 ( .INP(n2362), .ZN(n1109) );
  INVX0 U1249 ( .INP(n2362), .ZN(n1110) );
  MUX41X1 U1250 ( .IN1(\regf[16][13] ), .IN3(\regf[18][13] ), .IN2(
        \regf[17][13] ), .IN4(\regf[19][13] ), .S0(n1342), .S1(n1443), .Q(
        n1577) );
  MUX41X1 U1251 ( .IN1(\regf[12][31] ), .IN3(\regf[14][31] ), .IN2(
        \regf[13][31] ), .IN4(\regf[15][31] ), .S0(n1348), .S1(n1080), .Q(
        n1759) );
  MUX41X1 U1252 ( .IN1(\regf[12][30] ), .IN3(\regf[14][30] ), .IN2(
        \regf[13][30] ), .IN4(\regf[15][30] ), .S0(n1347), .S1(n1434), .Q(
        n1749) );
  DELLN1X2 U1253 ( .INP(n1425), .Z(n1111) );
  MUX41X1 U1254 ( .IN1(\regf[4][31] ), .IN3(\regf[6][31] ), .IN2(\regf[5][31] ), .IN4(\regf[7][31] ), .S0(n1343), .S1(n1196), .Q(n1761) );
  MUX41X1 U1255 ( .IN1(\regf[20][19] ), .IN3(\regf[22][19] ), .IN2(
        \regf[21][19] ), .IN4(\regf[23][19] ), .S0(n1352), .S1(n1196), .Q(
        n1636) );
  MUX41X1 U1256 ( .IN1(\regf[16][27] ), .IN3(\regf[18][27] ), .IN2(
        \regf[17][27] ), .IN4(\regf[19][27] ), .S0(n1352), .S1(n1175), .Q(
        n1717) );
  MUX41X1 U1257 ( .IN1(\regf[16][23] ), .IN3(\regf[18][23] ), .IN2(
        \regf[17][23] ), .IN4(\regf[19][23] ), .S0(n1348), .S1(n1120), .Q(
        n1677) );
  MUX41X1 U1258 ( .IN1(\regf[16][12] ), .IN3(\regf[18][12] ), .IN2(
        \regf[17][12] ), .IN4(\regf[19][12] ), .S0(n1343), .S1(n1158), .Q(
        n1567) );
  MUX41X1 U1259 ( .IN1(\regf[16][22] ), .IN3(\regf[18][22] ), .IN2(
        \regf[17][22] ), .IN4(\regf[19][22] ), .S0(n1347), .S1(n1151), .Q(
        n1667) );
  DELLN1X2 U1260 ( .INP(n1388), .Z(n1112) );
  MUX41X2 U1261 ( .IN1(n2064), .IN3(n2062), .IN2(n2063), .IN4(n2061), .S0(
        n2377), .S1(n2371), .Q(n2065) );
  NAND3X1 U1262 ( .IN1(\regf[3][2] ), .IN2(n1284), .IN3(n1132), .QN(n1882) );
  INVX0 U1263 ( .INP(n1369), .ZN(n1113) );
  NAND3X1 U1264 ( .IN1(\regf[3][23] ), .IN2(n1291), .IN3(n1438), .QN(n1798) );
  MUX21X2 U1265 ( .IN1(n2070), .IN2(n2065), .S(n2381), .Q(rd_dataB[15]) );
  MUX41X1 U1266 ( .IN1(\regf[4][21] ), .IN3(\regf[6][21] ), .IN2(\regf[5][21] ), .IN4(\regf[7][21] ), .S0(n1345), .S1(n1194), .Q(n1661) );
  MUX41X1 U1267 ( .IN1(\regf[16][30] ), .IN3(\regf[18][30] ), .IN2(
        \regf[17][30] ), .IN4(\regf[19][30] ), .S0(n1342), .S1(n1194), .Q(
        n1747) );
  NAND3X1 U1268 ( .IN1(\regf[3][24] ), .IN2(n1205), .IN3(n1366), .QN(n2261) );
  NAND3X1 U1269 ( .IN1(\regf[3][11] ), .IN2(n1126), .IN3(n1106), .QN(n2313) );
  MUX41X2 U1270 ( .IN1(\regf[4][22] ), .IN3(\regf[6][22] ), .IN2(\regf[5][22] ), .IN4(\regf[7][22] ), .S0(n1347), .S1(n1123), .Q(n1671) );
  DELLN1X2 U1271 ( .INP(n1424), .Z(n1114) );
  DELLN1X2 U1272 ( .INP(n1424), .Z(n1115) );
  INVX0 U1273 ( .INP(n1370), .ZN(n1116) );
  MUX41X1 U1274 ( .IN1(\regf[17][17] ), .IN3(\regf[19][17] ), .IN2(
        \regf[16][17] ), .IN4(\regf[18][17] ), .S0(n1233), .S1(n2364), .Q(
        n2084) );
  DELLN1X2 U1275 ( .INP(n1892), .Z(n1894) );
  NAND3X1 U1276 ( .IN1(\regf[3][15] ), .IN2(n1295), .IN3(n1195), .QN(n1830) );
  NAND3X1 U1277 ( .IN1(\regf[3][30] ), .IN2(n1287), .IN3(n1195), .QN(n1770) );
  NAND3X1 U1278 ( .IN1(\regf[3][24] ), .IN2(n1284), .IN3(n1183), .QN(n1794) );
  DELLN1X2 U1279 ( .INP(n1369), .Z(n2364) );
  INVX0 U1280 ( .INP(n1243), .ZN(n1117) );
  OR2X1 U1281 ( .IN1(n1118), .IN2(n1422), .Q(n1865) );
  INVX0 U1282 ( .INP(n1894), .ZN(n1119) );
  MUX21X2 U1283 ( .IN1(n1884), .IN2(n1885), .S(n1309), .Q(n1887) );
  DELLN1X2 U1284 ( .INP(n1426), .Z(n1120) );
  DELLN1X2 U1285 ( .INP(n1426), .Z(n1121) );
  OR2X1 U1286 ( .IN1(n1122), .IN2(n1395), .Q(n2308) );
  MUX41X1 U1287 ( .IN1(\regf[25][12] ), .IN3(\regf[27][12] ), .IN2(
        \regf[24][12] ), .IN4(\regf[26][12] ), .S0(n1287), .S1(n1894), .Q(
        n1565) );
  DELLN1X2 U1288 ( .INP(n1424), .Z(n1123) );
  DELLN1X2 U1289 ( .INP(n1417), .Z(n1124) );
  MUX41X1 U1290 ( .IN1(\regf[25][23] ), .IN3(\regf[27][23] ), .IN2(
        \regf[24][23] ), .IN4(\regf[26][23] ), .S0(n1292), .S1(n1403), .Q(
        n1675) );
  INVX0 U1291 ( .INP(n1239), .ZN(n1125) );
  INVX0 U1292 ( .INP(n1239), .ZN(n1126) );
  DELLN1X2 U1293 ( .INP(n1425), .Z(n1127) );
  DELLN1X2 U1294 ( .INP(n1425), .Z(n1128) );
  DELLN1X2 U1295 ( .INP(n1424), .Z(n1129) );
  INVX0 U1296 ( .INP(n2363), .ZN(n1130) );
  DELLN1X2 U1297 ( .INP(n1368), .Z(n2361) );
  MUX41X1 U1298 ( .IN1(\regf[5][27] ), .IN3(\regf[7][27] ), .IN2(\regf[4][27] ), .IN4(\regf[6][27] ), .S0(n1352), .S1(n1083), .Q(n1721) );
  DELLN1X2 U1299 ( .INP(n1416), .Z(n1131) );
  DELLN1X2 U1300 ( .INP(n1416), .Z(n1132) );
  INVX0 U1301 ( .INP(n2361), .ZN(n1133) );
  INVX0 U1302 ( .INP(n1279), .ZN(n1134) );
  DELLN1X2 U1303 ( .INP(n1380), .Z(n1135) );
  DELLN1X2 U1304 ( .INP(n1380), .Z(n1182) );
  OR2X1 U1305 ( .IN1(n1136), .IN2(n1389), .Q(n2300) );
  MUX21X2 U1306 ( .IN1(n1796), .IN2(n1797), .S(n1296), .Q(n1799) );
  DELLN1X2 U1307 ( .INP(n1425), .Z(n1180) );
  INVX0 U1308 ( .INP(n1369), .ZN(n1137) );
  INVX0 U1309 ( .INP(n2361), .ZN(n1138) );
  INVX0 U1310 ( .INP(n2361), .ZN(n1139) );
  DELLN1X2 U1311 ( .INP(n1379), .Z(n1140) );
  DELLN1X2 U1312 ( .INP(n1388), .Z(n1141) );
  DELLN1X2 U1313 ( .INP(n1424), .Z(n1174) );
  DELLN1X2 U1314 ( .INP(n1379), .Z(n1142) );
  DELLN1X2 U1315 ( .INP(n1388), .Z(n1143) );
  NAND3X1 U1316 ( .IN1(\regf[3][25] ), .IN2(n1328), .IN3(n1175), .QN(n1790) );
  NAND3X1 U1317 ( .IN1(\regf[3][8] ), .IN2(n1328), .IN3(n1432), .QN(n1858) );
  DELLN1X2 U1318 ( .INP(n1424), .Z(n1185) );
  DELLN1X2 U1319 ( .INP(n1371), .Z(n1165) );
  OR2X1 U1320 ( .IN1(n1144), .IN2(n1422), .Q(n1801) );
  NAND3X1 U1321 ( .IN1(\regf[3][4] ), .IN2(n1300), .IN3(n1397), .QN(n1874) );
  DELLN1X2 U1322 ( .INP(n1426), .Z(n1177) );
  DELLN1X2 U1323 ( .INP(n1417), .Z(n1183) );
  MUX41X1 U1324 ( .IN1(\regf[25][23] ), .IN3(\regf[27][23] ), .IN2(
        \regf[24][23] ), .IN4(\regf[26][23] ), .S0(n1213), .S1(n2364), .Q(
        n2142) );
  DELLN1X2 U1325 ( .INP(n2360), .Z(n2363) );
  NAND3X1 U1326 ( .IN1(\regf[3][4] ), .IN2(n1263), .IN3(n1389), .QN(n2341) );
  NAND3X1 U1327 ( .IN1(\regf[3][26] ), .IN2(n1215), .IN3(n1354), .QN(n2253) );
  MUX21X2 U1328 ( .IN1(n2303), .IN2(n2304), .S(n1233), .Q(n2306) );
  MUX21X2 U1329 ( .IN1(n2231), .IN2(n2232), .S(n1212), .Q(n2234) );
  MUX21X2 U1330 ( .IN1(n2239), .IN2(n2240), .S(n1213), .Q(n2242) );
  DELLN1X2 U1331 ( .INP(n1426), .Z(n1172) );
  MUX21X2 U1332 ( .IN1(n2347), .IN2(n2348), .S(n1228), .Q(n2350) );
  INVX0 U1333 ( .INP(n1369), .ZN(n1145) );
  MUX41X1 U1334 ( .IN1(\regf[25][25] ), .IN3(\regf[27][25] ), .IN2(
        \regf[24][25] ), .IN4(\regf[26][25] ), .S0(n1215), .S1(n1356), .Q(
        n2162) );
  DELLN1X2 U1335 ( .INP(n1426), .Z(n1175) );
  DELLN1X2 U1336 ( .INP(n1416), .Z(n1194) );
  DELLN1X2 U1337 ( .INP(n1380), .Z(n1171) );
  DELLN1X2 U1338 ( .INP(n1380), .Z(n1181) );
  DELLN1X2 U1339 ( .INP(n1417), .Z(n1197) );
  DELLN1X2 U1340 ( .INP(n1425), .Z(n1178) );
  DELLN1X2 U1341 ( .INP(n1371), .Z(n1163) );
  DELLN1X2 U1342 ( .INP(n1378), .Z(n1169) );
  DELLN1X2 U1343 ( .INP(n1380), .Z(n1168) );
  DELLN1X2 U1344 ( .INP(n1103), .Z(n1166) );
  DELLN1X2 U1345 ( .INP(n1379), .Z(n1188) );
  NAND3X1 U1346 ( .IN1(\regf[3][23] ), .IN2(n1257), .IN3(n1376), .QN(n2265) );
  NAND3X1 U1347 ( .IN1(\regf[3][21] ), .IN2(n1335), .IN3(n1084), .QN(n1806) );
  NAND3X1 U1348 ( .IN1(\regf[3][22] ), .IN2(n1301), .IN3(n1436), .QN(n1802) );
  NAND3X1 U1349 ( .IN1(\regf[3][20] ), .IN2(n1335), .IN3(n1438), .QN(n1810) );
  NAND3X1 U1350 ( .IN1(\regf[3][17] ), .IN2(n1335), .IN3(n1443), .QN(n1822) );
  NAND3X1 U1351 ( .IN1(\regf[3][19] ), .IN2(n1335), .IN3(n1085), .QN(n1814) );
  NAND3X1 U1352 ( .IN1(\regf[3][21] ), .IN2(n1207), .IN3(n1116), .QN(n2273) );
  NAND3X1 U1353 ( .IN1(\regf[3][22] ), .IN2(n1258), .IN3(n1396), .QN(n2269) );
  NAND3X1 U1354 ( .IN1(\regf[3][20] ), .IN2(n1256), .IN3(n1357), .QN(n2277) );
  NAND3X1 U1355 ( .IN1(\regf[3][17] ), .IN2(n1254), .IN3(n1186), .QN(n2289) );
  NAND3X1 U1356 ( .IN1(\regf[3][19] ), .IN2(n1255), .IN3(n1363), .QN(n2281) );
  NAND3X1 U1357 ( .IN1(\regf[3][0] ), .IN2(n1218), .IN3(n1394), .QN(n2357) );
  DELLN1X2 U1358 ( .INP(n1379), .Z(n1191) );
  INVX0 U1359 ( .INP(n1414), .ZN(n1146) );
  NAND3X1 U1360 ( .IN1(\regf[3][27] ), .IN2(n1214), .IN3(n1113), .QN(n2249) );
  NAND3X1 U1361 ( .IN1(\regf[3][27] ), .IN2(n1285), .IN3(n1429), .QN(n1782) );
  NAND3X1 U1362 ( .IN1(\regf[3][12] ), .IN2(n1251), .IN3(n1354), .QN(n2309) );
  NAND3X1 U1363 ( .IN1(\regf[3][7] ), .IN2(n1245), .IN3(n1386), .QN(n2329) );
  NAND3X1 U1364 ( .IN1(\regf[3][9] ), .IN2(n1252), .IN3(n1187), .QN(n2321) );
  NAND3X1 U1365 ( .IN1(\regf[3][5] ), .IN2(n1261), .IN3(n1386), .QN(n2337) );
  NAND3X1 U1366 ( .IN1(\regf[3][28] ), .IN2(n1213), .IN3(n1386), .QN(n2245) );
  NAND3X1 U1367 ( .IN1(\regf[3][12] ), .IN2(n1299), .IN3(n1436), .QN(n1842) );
  NAND3X1 U1368 ( .IN1(\regf[3][7] ), .IN2(n1327), .IN3(n1433), .QN(n1862) );
  NAND3X1 U1369 ( .IN1(\regf[3][9] ), .IN2(n1333), .IN3(n1431), .QN(n1854) );
  NAND3X1 U1370 ( .IN1(\regf[3][5] ), .IN2(n1134), .IN3(n1075), .QN(n1870) );
  NAND3X1 U1371 ( .IN1(\regf[3][28] ), .IN2(n1293), .IN3(n1076), .QN(n1778) );
  NAND3X1 U1372 ( .IN1(\regf[3][3] ), .IN2(n1217), .IN3(n1386), .QN(n2345) );
  NAND3X1 U1373 ( .IN1(\regf[3][3] ), .IN2(n1298), .IN3(n1437), .QN(n1878) );
  DELLN1X2 U1374 ( .INP(n1373), .Z(n1147) );
  DELLN1X2 U1375 ( .INP(n1373), .Z(n1148) );
  DELLN1X2 U1376 ( .INP(n1425), .Z(n1149) );
  DELLN1X2 U1377 ( .INP(n1442), .Z(n1150) );
  DELLN1X2 U1378 ( .INP(n1400), .Z(n1151) );
  DELLN1X2 U1379 ( .INP(n1373), .Z(n1152) );
  DELLN1X2 U1380 ( .INP(n1388), .Z(n1153) );
  DELLN1X2 U1381 ( .INP(n1379), .Z(n1154) );
  DELLN1X2 U1382 ( .INP(n1371), .Z(n1155) );
  DELLN1X2 U1383 ( .INP(n1103), .Z(n1156) );
  DELLN1X2 U1384 ( .INP(n1379), .Z(n1157) );
  DELLN1X2 U1385 ( .INP(n1420), .Z(n1158) );
  DELLN1X2 U1386 ( .INP(n1417), .Z(n1159) );
  DELLN1X2 U1387 ( .INP(n1420), .Z(n1160) );
  DELLN1X2 U1388 ( .INP(n1416), .Z(n1161) );
  DELLN1X2 U1389 ( .INP(n1420), .Z(n1162) );
  NAND3X1 U1390 ( .IN1(\regf[3][14] ), .IN2(n1247), .IN3(n1366), .QN(n2301) );
  NAND3X1 U1391 ( .IN1(\regf[3][18] ), .IN2(n1247), .IN3(n1147), .QN(n2285) );
  NAND3X1 U1392 ( .IN1(\regf[3][14] ), .IN2(n1327), .IN3(n1159), .QN(n1834) );
  NAND3X1 U1393 ( .IN1(\regf[3][18] ), .IN2(n1297), .IN3(n1435), .QN(n1818) );
  DELLN1X2 U1394 ( .INP(n1378), .Z(n1164) );
  DELLN1X2 U1395 ( .INP(n1380), .Z(n1167) );
  DELLN1X2 U1396 ( .INP(n1388), .Z(n1170) );
  DELLN1X2 U1397 ( .INP(n1425), .Z(n1173) );
  DELLN1X2 U1398 ( .INP(n1426), .Z(n1176) );
  DELLN1X2 U1399 ( .INP(n1425), .Z(n1179) );
  DELLN1X2 U1400 ( .INP(n1424), .Z(n1184) );
  DELLN1X2 U1401 ( .INP(n1103), .Z(n1189) );
  DELLN1X2 U1402 ( .INP(n1375), .Z(n1186) );
  DELLN1X2 U1403 ( .INP(n1420), .Z(n1195) );
  DELLN1X2 U1404 ( .INP(n1420), .Z(n1192) );
  DELLN1X2 U1405 ( .INP(n1378), .Z(n1187) );
  DELLN1X2 U1406 ( .INP(n1378), .Z(n1190) );
  DELLN1X2 U1407 ( .INP(n1416), .Z(n1193) );
  DELLN1X2 U1408 ( .INP(n1417), .Z(n1196) );
  INVX0 U1409 ( .INP(N17), .ZN(n1198) );
  INVX0 U1410 ( .INP(N17), .ZN(n1199) );
  INVX0 U1411 ( .INP(N17), .ZN(n1200) );
  INVX0 U1412 ( .INP(N17), .ZN(n1201) );
  INVX0 U1413 ( .INP(N17), .ZN(n1202) );
  INVX0 U1414 ( .INP(N17), .ZN(n1203) );
  INVX0 U1415 ( .INP(n1198), .ZN(n1204) );
  INVX0 U1416 ( .INP(n1198), .ZN(n1205) );
  INVX0 U1417 ( .INP(n1198), .ZN(n1206) );
  INVX0 U1418 ( .INP(n1198), .ZN(n1207) );
  INVX0 U1419 ( .INP(n1198), .ZN(n1208) );
  INVX0 U1420 ( .INP(n1199), .ZN(n1209) );
  INVX0 U1421 ( .INP(n1199), .ZN(n1210) );
  INVX0 U1422 ( .INP(n1199), .ZN(n1211) );
  INVX0 U1423 ( .INP(n1199), .ZN(n1212) );
  INVX0 U1424 ( .INP(n1199), .ZN(n1213) );
  INVX0 U1425 ( .INP(n1201), .ZN(n1214) );
  INVX0 U1426 ( .INP(n1202), .ZN(n1215) );
  INVX0 U1427 ( .INP(n1199), .ZN(n1216) );
  INVX0 U1428 ( .INP(n1198), .ZN(n1217) );
  INVX0 U1429 ( .INP(n1200), .ZN(n1218) );
  INVX0 U1430 ( .INP(n1200), .ZN(n1219) );
  INVX0 U1431 ( .INP(n1200), .ZN(n1220) );
  INVX0 U1432 ( .INP(n1200), .ZN(n1221) );
  INVX0 U1433 ( .INP(n1200), .ZN(n1222) );
  INVX0 U1434 ( .INP(n1200), .ZN(n1223) );
  INVX0 U1435 ( .INP(n1201), .ZN(n1224) );
  INVX0 U1436 ( .INP(n1201), .ZN(n1225) );
  INVX0 U1437 ( .INP(n1201), .ZN(n1226) );
  INVX0 U1438 ( .INP(n1201), .ZN(n1227) );
  INVX0 U1439 ( .INP(n1201), .ZN(n1228) );
  INVX0 U1440 ( .INP(n1202), .ZN(n1229) );
  INVX0 U1441 ( .INP(n1200), .ZN(n1230) );
  INVX0 U1442 ( .INP(n1201), .ZN(n1231) );
  INVX0 U1443 ( .INP(n1202), .ZN(n1232) );
  INVX0 U1444 ( .INP(n1202), .ZN(n1233) );
  INVX0 U1445 ( .INP(n1202), .ZN(n1234) );
  INVX0 U1446 ( .INP(n1202), .ZN(n1235) );
  INVX0 U1447 ( .INP(n1203), .ZN(n1236) );
  INVX0 U1448 ( .INP(n1203), .ZN(n1237) );
  INVX0 U1449 ( .INP(n1203), .ZN(n1238) );
  INVX0 U1450 ( .INP(n2367), .ZN(n1239) );
  INVX0 U1451 ( .INP(n2367), .ZN(n1240) );
  INVX0 U1452 ( .INP(n2367), .ZN(n1241) );
  INVX0 U1453 ( .INP(n2367), .ZN(n1242) );
  INVX0 U1454 ( .INP(n2367), .ZN(n1243) );
  INVX0 U1455 ( .INP(n2367), .ZN(n1244) );
  INVX0 U1456 ( .INP(n1239), .ZN(n1245) );
  INVX0 U1457 ( .INP(n1239), .ZN(n1246) );
  INVX0 U1458 ( .INP(n1239), .ZN(n1247) );
  INVX0 U1459 ( .INP(n1240), .ZN(n1248) );
  INVX0 U1460 ( .INP(n1240), .ZN(n1249) );
  INVX0 U1461 ( .INP(n1240), .ZN(n1250) );
  INVX0 U1462 ( .INP(n1240), .ZN(n1251) );
  INVX0 U1463 ( .INP(n1240), .ZN(n1252) );
  INVX0 U1464 ( .INP(n1241), .ZN(n1253) );
  INVX0 U1465 ( .INP(n1241), .ZN(n1254) );
  INVX0 U1466 ( .INP(n1241), .ZN(n1255) );
  INVX0 U1467 ( .INP(n1241), .ZN(n1256) );
  INVX0 U1468 ( .INP(n1242), .ZN(n1257) );
  INVX0 U1469 ( .INP(n1242), .ZN(n1258) );
  INVX0 U1470 ( .INP(n1242), .ZN(n1259) );
  INVX0 U1471 ( .INP(n1242), .ZN(n1260) );
  INVX0 U1472 ( .INP(n1243), .ZN(n1261) );
  INVX0 U1473 ( .INP(n1243), .ZN(n1262) );
  INVX0 U1474 ( .INP(n1243), .ZN(n1263) );
  INVX0 U1475 ( .INP(n1243), .ZN(n1264) );
  INVX0 U1476 ( .INP(n1203), .ZN(n1265) );
  INVX0 U1477 ( .INP(n1203), .ZN(n1266) );
  INVX0 U1478 ( .INP(n1203), .ZN(n1267) );
  INVX0 U1479 ( .INP(n1241), .ZN(n1268) );
  INVX0 U1480 ( .INP(n1242), .ZN(n1269) );
  INVX0 U1481 ( .INP(n1239), .ZN(n1270) );
  INVX0 U1482 ( .INP(n1244), .ZN(n1271) );
  INVX0 U1483 ( .INP(n1244), .ZN(n1272) );
  INVX0 U1484 ( .INP(n1244), .ZN(n1273) );
  INVX0 U1485 ( .INP(n1244), .ZN(n1274) );
  INVX0 U1486 ( .INP(n1244), .ZN(n1275) );
  INVX0 U1487 ( .INP(N12), .ZN(n1276) );
  INVX0 U1488 ( .INP(N12), .ZN(n1277) );
  INVX0 U1489 ( .INP(N12), .ZN(n1278) );
  INVX0 U1490 ( .INP(N12), .ZN(n1279) );
  INVX0 U1491 ( .INP(N12), .ZN(n1280) );
  INVX0 U1492 ( .INP(N12), .ZN(n1281) );
  INVX0 U1493 ( .INP(N12), .ZN(n1282) );
  INVX0 U1494 ( .INP(n1276), .ZN(n1283) );
  INVX0 U1495 ( .INP(n1276), .ZN(n1284) );
  INVX0 U1496 ( .INP(n1276), .ZN(n1285) );
  INVX0 U1497 ( .INP(n1276), .ZN(n1286) );
  INVX0 U1498 ( .INP(n1276), .ZN(n1287) );
  INVX0 U1499 ( .INP(n1276), .ZN(n1288) );
  INVX0 U1500 ( .INP(n1276), .ZN(n1289) );
  INVX0 U1501 ( .INP(n1281), .ZN(n1290) );
  INVX0 U1502 ( .INP(n1280), .ZN(n1291) );
  INVX0 U1503 ( .INP(n1282), .ZN(n1292) );
  INVX0 U1504 ( .INP(n1277), .ZN(n1293) );
  INVX0 U1505 ( .INP(n1277), .ZN(n1294) );
  INVX0 U1506 ( .INP(n1277), .ZN(n1295) );
  INVX0 U1507 ( .INP(n1277), .ZN(n1296) );
  INVX0 U1508 ( .INP(n1277), .ZN(n1297) );
  INVX0 U1509 ( .INP(n1278), .ZN(n1298) );
  INVX0 U1510 ( .INP(n1278), .ZN(n1299) );
  INVX0 U1511 ( .INP(n1278), .ZN(n1300) );
  INVX0 U1512 ( .INP(n1278), .ZN(n1301) );
  INVX0 U1513 ( .INP(n1278), .ZN(n1302) );
  INVX0 U1514 ( .INP(n1279), .ZN(n1303) );
  INVX0 U1515 ( .INP(n1279), .ZN(n1304) );
  INVX0 U1516 ( .INP(n1279), .ZN(n1305) );
  INVX0 U1517 ( .INP(n1279), .ZN(n1306) );
  INVX0 U1518 ( .INP(n1279), .ZN(n1307) );
  INVX0 U1519 ( .INP(n1280), .ZN(n1308) );
  INVX0 U1520 ( .INP(n1280), .ZN(n1309) );
  INVX0 U1521 ( .INP(n1280), .ZN(n1310) );
  INVX0 U1522 ( .INP(n1281), .ZN(n1311) );
  INVX0 U1523 ( .INP(n1281), .ZN(n1312) );
  INVX0 U1524 ( .INP(n1281), .ZN(n1313) );
  INVX0 U1525 ( .INP(n1281), .ZN(n1314) );
  INVX0 U1526 ( .INP(n1282), .ZN(n1315) );
  INVX0 U1527 ( .INP(n1282), .ZN(n1316) );
  INVX0 U1528 ( .INP(n1282), .ZN(n1317) );
  INVX0 U1529 ( .INP(n1282), .ZN(n1318) );
  INVX0 U1530 ( .INP(n1282), .ZN(n1319) );
  INVX0 U1531 ( .INP(n1895), .ZN(n1320) );
  INVX0 U1532 ( .INP(n1895), .ZN(n1321) );
  INVX0 U1533 ( .INP(n1895), .ZN(n1322) );
  INVX0 U1534 ( .INP(n1895), .ZN(n1323) );
  INVX0 U1535 ( .INP(n1895), .ZN(n1324) );
  INVX0 U1536 ( .INP(n1322), .ZN(n1325) );
  INVX0 U1537 ( .INP(n1323), .ZN(n1326) );
  INVX0 U1538 ( .INP(n1324), .ZN(n1327) );
  INVX0 U1539 ( .INP(n1324), .ZN(n1328) );
  INVX0 U1540 ( .INP(n1321), .ZN(n1329) );
  INVX0 U1541 ( .INP(n1324), .ZN(n1330) );
  INVX0 U1542 ( .INP(n1320), .ZN(n1331) );
  INVX0 U1543 ( .INP(n1323), .ZN(n1332) );
  INVX0 U1544 ( .INP(n1279), .ZN(n1333) );
  INVX0 U1545 ( .INP(n1279), .ZN(n1334) );
  INVX0 U1546 ( .INP(n1320), .ZN(n1335) );
  INVX0 U1547 ( .INP(n1321), .ZN(n1336) );
  INVX0 U1548 ( .INP(n1321), .ZN(n1337) );
  INVX0 U1549 ( .INP(n1324), .ZN(n1338) );
  INVX0 U1550 ( .INP(n1323), .ZN(n1339) );
  INVX0 U1551 ( .INP(n1320), .ZN(n1340) );
  INVX0 U1552 ( .INP(n1322), .ZN(n1341) );
  INVX0 U1553 ( .INP(n1323), .ZN(n1342) );
  INVX0 U1554 ( .INP(n1320), .ZN(n1343) );
  INVX0 U1555 ( .INP(n1322), .ZN(n1344) );
  INVX0 U1556 ( .INP(n1276), .ZN(n1345) );
  INVX0 U1557 ( .INP(n1281), .ZN(n1346) );
  INVX0 U1558 ( .INP(n1323), .ZN(n1347) );
  INVX0 U1559 ( .INP(n1280), .ZN(n1348) );
  INVX0 U1560 ( .INP(n1320), .ZN(n1349) );
  INVX0 U1561 ( .INP(n1321), .ZN(n1350) );
  INVX0 U1562 ( .INP(n1322), .ZN(n1351) );
  INVX0 U1563 ( .INP(n1321), .ZN(n1352) );
  INVX0 U1564 ( .INP(n1322), .ZN(n1353) );
  INVX0 U1565 ( .INP(n2360), .ZN(n1354) );
  INVX0 U1566 ( .INP(n2359), .ZN(n1355) );
  INVX0 U1567 ( .INP(n1389), .ZN(n1356) );
  INVX0 U1568 ( .INP(n2362), .ZN(n1357) );
  INVX0 U1569 ( .INP(n2363), .ZN(n1358) );
  INVX0 U1570 ( .INP(n2361), .ZN(n1359) );
  INVX0 U1571 ( .INP(n1373), .ZN(n1360) );
  INVX0 U1572 ( .INP(n1373), .ZN(n1361) );
  INVX0 U1573 ( .INP(n2366), .ZN(n1362) );
  INVX0 U1574 ( .INP(n1370), .ZN(n1363) );
  INVX0 U1575 ( .INP(n2359), .ZN(n1364) );
  INVX0 U1576 ( .INP(n2365), .ZN(n1365) );
  INVX0 U1577 ( .INP(n1370), .ZN(n1366) );
  INVX0 U1578 ( .INP(N16), .ZN(n1367) );
  INVX0 U1579 ( .INP(N16), .ZN(n1368) );
  INVX0 U1580 ( .INP(N16), .ZN(n1369) );
  INVX0 U1581 ( .INP(N16), .ZN(n1370) );
  INVX0 U1582 ( .INP(n1368), .ZN(n1371) );
  INVX0 U1583 ( .INP(n1367), .ZN(n1372) );
  INVX0 U1584 ( .INP(n2359), .ZN(n1373) );
  INVX0 U1585 ( .INP(n2360), .ZN(n1374) );
  INVX0 U1586 ( .INP(n1367), .ZN(n1375) );
  INVX0 U1587 ( .INP(n2359), .ZN(n1376) );
  INVX0 U1588 ( .INP(n1370), .ZN(n1377) );
  INVX0 U1589 ( .INP(n1368), .ZN(n1378) );
  INVX0 U1590 ( .INP(n1367), .ZN(n1379) );
  INVX0 U1591 ( .INP(n1368), .ZN(n1380) );
  INVX0 U1592 ( .INP(n2359), .ZN(n1381) );
  INVX0 U1593 ( .INP(n2359), .ZN(n1382) );
  INVX0 U1594 ( .INP(n1369), .ZN(n1383) );
  INVX0 U1595 ( .INP(n1370), .ZN(n1384) );
  INVX0 U1596 ( .INP(n1369), .ZN(n1385) );
  INVX0 U1597 ( .INP(n1369), .ZN(n1386) );
  INVX0 U1598 ( .INP(n1369), .ZN(n1387) );
  INVX0 U1599 ( .INP(n1367), .ZN(n1388) );
  INVX0 U1600 ( .INP(n1368), .ZN(n1389) );
  INVX0 U1601 ( .INP(n1370), .ZN(n1390) );
  INVX0 U1602 ( .INP(n1367), .ZN(n1391) );
  INVX0 U1603 ( .INP(n1367), .ZN(n1392) );
  INVX0 U1604 ( .INP(n1370), .ZN(n1393) );
  INVX0 U1605 ( .INP(n1370), .ZN(n1394) );
  INVX0 U1606 ( .INP(n1369), .ZN(n1395) );
  INVX0 U1607 ( .INP(n1370), .ZN(n1396) );
  DELLN1X2 U1608 ( .INP(n2360), .Z(n2365) );
  DELLN1X2 U1609 ( .INP(n2360), .Z(n2366) );
  INVX0 U1610 ( .INP(n1412), .ZN(n1397) );
  INVX0 U1611 ( .INP(n1411), .ZN(n1398) );
  INVX0 U1612 ( .INP(n1398), .ZN(n1399) );
  INVX0 U1613 ( .INP(n1414), .ZN(n1400) );
  INVX0 U1614 ( .INP(n1397), .ZN(n1401) );
  INVX0 U1615 ( .INP(n1894), .ZN(n1402) );
  INVX0 U1616 ( .INP(n1442), .ZN(n1403) );
  INVX0 U1617 ( .INP(n1894), .ZN(n1404) );
  INVX0 U1618 ( .INP(n1415), .ZN(n1405) );
  INVX0 U1619 ( .INP(n1442), .ZN(n1406) );
  INVX0 U1620 ( .INP(n1894), .ZN(n1407) );
  INVX0 U1621 ( .INP(n1421), .ZN(n1408) );
  INVX0 U1622 ( .INP(n1415), .ZN(n1409) );
  INVX0 U1623 ( .INP(n1413), .ZN(n1410) );
  INVX0 U1624 ( .INP(N11), .ZN(n1411) );
  INVX0 U1625 ( .INP(N11), .ZN(n1412) );
  INVX0 U1626 ( .INP(N11), .ZN(n1413) );
  INVX0 U1627 ( .INP(N11), .ZN(n1414) );
  INVX0 U1628 ( .INP(N11), .ZN(n1415) );
  INVX0 U1629 ( .INP(n1411), .ZN(n1416) );
  INVX0 U1630 ( .INP(n1892), .ZN(n1417) );
  INVX0 U1631 ( .INP(n1412), .ZN(n1418) );
  INVX0 U1632 ( .INP(n1412), .ZN(n1419) );
  INVX0 U1633 ( .INP(n1892), .ZN(n1420) );
  INVX0 U1634 ( .INP(n1411), .ZN(n1421) );
  INVX0 U1635 ( .INP(n1413), .ZN(n1422) );
  INVX0 U1636 ( .INP(n1412), .ZN(n1423) );
  INVX0 U1637 ( .INP(n1411), .ZN(n1424) );
  INVX0 U1638 ( .INP(n1892), .ZN(n1425) );
  INVX0 U1639 ( .INP(n1412), .ZN(n1426) );
  INVX0 U1640 ( .INP(n1412), .ZN(n1427) );
  INVX0 U1641 ( .INP(n1413), .ZN(n1428) );
  INVX0 U1642 ( .INP(n1413), .ZN(n1429) );
  INVX0 U1643 ( .INP(n1415), .ZN(n1430) );
  INVX0 U1644 ( .INP(n1413), .ZN(n1431) );
  INVX0 U1645 ( .INP(n1413), .ZN(n1432) );
  INVX0 U1646 ( .INP(n1413), .ZN(n1433) );
  INVX0 U1647 ( .INP(n1414), .ZN(n1434) );
  INVX0 U1648 ( .INP(n1414), .ZN(n1435) );
  INVX0 U1649 ( .INP(n1414), .ZN(n1436) );
  INVX0 U1650 ( .INP(n1414), .ZN(n1437) );
  INVX0 U1651 ( .INP(n1414), .ZN(n1438) );
  INVX0 U1652 ( .INP(n1415), .ZN(n1439) );
  INVX0 U1653 ( .INP(n1415), .ZN(n1440) );
  INVX0 U1654 ( .INP(n1415), .ZN(n1441) );
  INVX0 U1655 ( .INP(n1411), .ZN(n1442) );
  INVX0 U1656 ( .INP(n1415), .ZN(n1443) );
  DELLN1X2 U1657 ( .INP(n1368), .Z(n2362) );
  INVX0 U1658 ( .INP(n37), .ZN(n2523) );
  INVX0 U1659 ( .INP(n37), .ZN(n2524) );
  INVX0 U1660 ( .INP(n40), .ZN(n2518) );
  INVX0 U1661 ( .INP(n40), .ZN(n2519) );
  INVX0 U1662 ( .INP(n42), .ZN(n2513) );
  INVX0 U1663 ( .INP(n42), .ZN(n2514) );
  INVX0 U1664 ( .INP(n55), .ZN(n2483) );
  INVX0 U1665 ( .INP(n55), .ZN(n2484) );
  INVX0 U1666 ( .INP(n73), .ZN(n2408) );
  INVX0 U1667 ( .INP(n73), .ZN(n2409) );
  INVX0 U1668 ( .INP(n54), .ZN(n2488) );
  INVX0 U1669 ( .INP(n54), .ZN(n2489) );
  INVX0 U1670 ( .INP(n72), .ZN(n2413) );
  INVX0 U1671 ( .INP(n72), .ZN(n2414) );
  INVX0 U1672 ( .INP(n56), .ZN(n2478) );
  INVX0 U1673 ( .INP(n56), .ZN(n2479) );
  INVX0 U1674 ( .INP(n74), .ZN(n2403) );
  INVX0 U1675 ( .INP(n74), .ZN(n2404) );
  INVX0 U1676 ( .INP(n44), .ZN(n2508) );
  INVX0 U1677 ( .INP(n44), .ZN(n2509) );
  INVX0 U1678 ( .INP(n46), .ZN(n2504) );
  INVX0 U1679 ( .INP(n46), .ZN(n2505) );
  INVX0 U1680 ( .INP(n48), .ZN(n2500) );
  INVX0 U1681 ( .INP(n48), .ZN(n2501) );
  INVX0 U1682 ( .INP(n50), .ZN(n2496) );
  INVX0 U1683 ( .INP(n50), .ZN(n2497) );
  INVX0 U1684 ( .INP(n64), .ZN(n2446) );
  INVX0 U1685 ( .INP(n63), .ZN(n2451) );
  INVX0 U1686 ( .INP(n61), .ZN(n2456) );
  INVX0 U1687 ( .INP(n65), .ZN(n2441) );
  INVX0 U1688 ( .INP(n66), .ZN(n2436) );
  INVX0 U1689 ( .INP(n67), .ZN(n2431) );
  INVX0 U1690 ( .INP(n68), .ZN(n2426) );
  INVX0 U1691 ( .INP(n69), .ZN(n2421) );
  INVX0 U1692 ( .INP(n52), .ZN(n2492) );
  INVX0 U1693 ( .INP(n52), .ZN(n2493) );
  INVX0 U1694 ( .INP(n70), .ZN(n2417) );
  INVX0 U1695 ( .INP(n70), .ZN(n2418) );
  INVX0 U1696 ( .INP(n75), .ZN(n2398) );
  INVX0 U1697 ( .INP(n75), .ZN(n2399) );
  INVX0 U1698 ( .INP(n76), .ZN(n2394) );
  INVX0 U1699 ( .INP(n76), .ZN(n2395) );
  INVX0 U1700 ( .INP(n77), .ZN(n2390) );
  INVX0 U1701 ( .INP(n77), .ZN(n2391) );
  INVX0 U1702 ( .INP(n78), .ZN(n2386) );
  INVX0 U1703 ( .INP(n78), .ZN(n2387) );
  INVX0 U1704 ( .INP(n57), .ZN(n2473) );
  INVX0 U1705 ( .INP(n57), .ZN(n2474) );
  INVX0 U1706 ( .INP(n58), .ZN(n2469) );
  INVX0 U1707 ( .INP(n58), .ZN(n2470) );
  INVX0 U1708 ( .INP(n59), .ZN(n2465) );
  INVX0 U1709 ( .INP(n59), .ZN(n2466) );
  INVX0 U1710 ( .INP(n60), .ZN(n2461) );
  INVX0 U1711 ( .INP(n60), .ZN(n2462) );
  INVX0 U1712 ( .INP(n64), .ZN(n2447) );
  INVX0 U1713 ( .INP(n64), .ZN(n2448) );
  INVX0 U1714 ( .INP(n63), .ZN(n2452) );
  INVX0 U1715 ( .INP(n63), .ZN(n2453) );
  INVX0 U1716 ( .INP(n61), .ZN(n2457) );
  INVX0 U1717 ( .INP(n61), .ZN(n2458) );
  INVX0 U1718 ( .INP(n65), .ZN(n2442) );
  INVX0 U1719 ( .INP(n65), .ZN(n2443) );
  INVX0 U1720 ( .INP(n66), .ZN(n2437) );
  INVX0 U1721 ( .INP(n66), .ZN(n2438) );
  INVX0 U1722 ( .INP(n67), .ZN(n2432) );
  INVX0 U1723 ( .INP(n67), .ZN(n2433) );
  INVX0 U1724 ( .INP(n68), .ZN(n2427) );
  INVX0 U1725 ( .INP(n68), .ZN(n2428) );
  INVX0 U1726 ( .INP(n69), .ZN(n2422) );
  INVX0 U1727 ( .INP(n69), .ZN(n2423) );
  NBUFFX2 U1728 ( .INP(n2704), .Z(n2702) );
  NBUFFX2 U1729 ( .INP(n2704), .Z(n2701) );
  NBUFFX2 U1730 ( .INP(n2704), .Z(n2700) );
  NBUFFX2 U1731 ( .INP(n2704), .Z(n2699) );
  NBUFFX2 U1732 ( .INP(n2704), .Z(n2698) );
  NBUFFX2 U1733 ( .INP(n2704), .Z(n2697) );
  NBUFFX2 U1734 ( .INP(n2704), .Z(n2696) );
  NBUFFX2 U1735 ( .INP(n2704), .Z(n2695) );
  NBUFFX2 U1736 ( .INP(n2704), .Z(n2694) );
  NBUFFX2 U1737 ( .INP(n2704), .Z(n2693) );
  NBUFFX2 U1738 ( .INP(n2704), .Z(n2692) );
  NBUFFX2 U1739 ( .INP(n2705), .Z(n2691) );
  NBUFFX2 U1740 ( .INP(n2705), .Z(n2690) );
  NBUFFX2 U1741 ( .INP(n2705), .Z(n2689) );
  NBUFFX2 U1742 ( .INP(n2705), .Z(n2688) );
  NBUFFX2 U1743 ( .INP(n2705), .Z(n2687) );
  NBUFFX2 U1744 ( .INP(n2705), .Z(n2686) );
  NBUFFX2 U1745 ( .INP(n2705), .Z(n2685) );
  NBUFFX2 U1746 ( .INP(n2705), .Z(n2684) );
  NBUFFX2 U1747 ( .INP(n2705), .Z(n2683) );
  NBUFFX2 U1748 ( .INP(n2705), .Z(n2682) );
  NBUFFX2 U1749 ( .INP(n2705), .Z(n2681) );
  NBUFFX2 U1750 ( .INP(n2705), .Z(n2680) );
  NBUFFX2 U1751 ( .INP(n2706), .Z(n2679) );
  NBUFFX2 U1752 ( .INP(n2706), .Z(n2678) );
  NBUFFX2 U1753 ( .INP(n2706), .Z(n2677) );
  NBUFFX2 U1754 ( .INP(n2706), .Z(n2676) );
  NBUFFX2 U1755 ( .INP(n2706), .Z(n2675) );
  NBUFFX2 U1756 ( .INP(n2706), .Z(n2674) );
  NBUFFX2 U1757 ( .INP(n2706), .Z(n2673) );
  NBUFFX2 U1758 ( .INP(n2706), .Z(n2672) );
  NBUFFX2 U1759 ( .INP(n2706), .Z(n2671) );
  NBUFFX2 U1760 ( .INP(n2706), .Z(n2670) );
  NBUFFX2 U1761 ( .INP(n2706), .Z(n2669) );
  NBUFFX2 U1762 ( .INP(n2706), .Z(n2668) );
  NBUFFX2 U1763 ( .INP(n2707), .Z(n2667) );
  NBUFFX2 U1764 ( .INP(n2707), .Z(n2666) );
  NBUFFX2 U1765 ( .INP(n2707), .Z(n2665) );
  NBUFFX2 U1766 ( .INP(n2707), .Z(n2664) );
  NBUFFX2 U1767 ( .INP(n2707), .Z(n2663) );
  NBUFFX2 U1768 ( .INP(n2707), .Z(n2662) );
  NBUFFX2 U1769 ( .INP(n2707), .Z(n2661) );
  NBUFFX2 U1770 ( .INP(n2707), .Z(n2660) );
  NBUFFX2 U1771 ( .INP(n2707), .Z(n2659) );
  NBUFFX2 U1772 ( .INP(n2707), .Z(n2658) );
  NBUFFX2 U1773 ( .INP(n2707), .Z(n2657) );
  NBUFFX2 U1774 ( .INP(n2707), .Z(n2656) );
  NBUFFX2 U1775 ( .INP(n2708), .Z(n2655) );
  NBUFFX2 U1776 ( .INP(n2708), .Z(n2654) );
  NBUFFX2 U1777 ( .INP(n2708), .Z(n2653) );
  NBUFFX2 U1778 ( .INP(n2708), .Z(n2652) );
  NBUFFX2 U1779 ( .INP(n2708), .Z(n2651) );
  NBUFFX2 U1780 ( .INP(n2708), .Z(n2650) );
  NBUFFX2 U1781 ( .INP(n2708), .Z(n2649) );
  NBUFFX2 U1782 ( .INP(n2708), .Z(n2648) );
  NBUFFX2 U1783 ( .INP(n2708), .Z(n2647) );
  NBUFFX2 U1784 ( .INP(n2708), .Z(n2646) );
  NBUFFX2 U1785 ( .INP(n2708), .Z(n2645) );
  NBUFFX2 U1786 ( .INP(n2708), .Z(n2644) );
  NBUFFX2 U1787 ( .INP(n2709), .Z(n2643) );
  NBUFFX2 U1788 ( .INP(n2709), .Z(n2642) );
  NBUFFX2 U1789 ( .INP(n2709), .Z(n2641) );
  NBUFFX2 U1790 ( .INP(n2709), .Z(n2640) );
  NBUFFX2 U1791 ( .INP(n2709), .Z(n2639) );
  NBUFFX2 U1792 ( .INP(n2709), .Z(n2638) );
  NBUFFX2 U1793 ( .INP(n2709), .Z(n2637) );
  NBUFFX2 U1794 ( .INP(n2709), .Z(n2636) );
  NBUFFX2 U1795 ( .INP(n2709), .Z(n2635) );
  NBUFFX2 U1796 ( .INP(n2709), .Z(n2634) );
  NBUFFX2 U1797 ( .INP(n2709), .Z(n2633) );
  NBUFFX2 U1798 ( .INP(n2709), .Z(n2632) );
  NBUFFX2 U1799 ( .INP(n2710), .Z(n2631) );
  NBUFFX2 U1800 ( .INP(n2710), .Z(n2630) );
  NBUFFX2 U1801 ( .INP(n2710), .Z(n2629) );
  NBUFFX2 U1802 ( .INP(n2710), .Z(n2628) );
  NBUFFX2 U1803 ( .INP(n2710), .Z(n2627) );
  NBUFFX2 U1804 ( .INP(n2710), .Z(n2626) );
  NBUFFX2 U1805 ( .INP(n2710), .Z(n2625) );
  NBUFFX2 U1806 ( .INP(n2710), .Z(n2624) );
  NBUFFX2 U1807 ( .INP(n2710), .Z(n2623) );
  NBUFFX2 U1808 ( .INP(n2710), .Z(n2622) );
  NBUFFX2 U1809 ( .INP(n2710), .Z(n2621) );
  NBUFFX2 U1810 ( .INP(n2704), .Z(n2703) );
  NAND2X0 U1811 ( .IN1(n1386), .IN2(\regf[1][30] ), .QN(n2235) );
  NAND2X0 U1812 ( .IN1(n1422), .IN2(\regf[1][30] ), .QN(n1768) );
  NAND2X0 U1813 ( .IN1(n2238), .IN2(n2237), .QN(n2219) );
  NAND2X0 U1814 ( .IN1(\regf[2][30] ), .IN2(n1360), .QN(n2236) );
  NAND2X0 U1815 ( .IN1(n1771), .IN2(n1770), .QN(n1752) );
  NAND2X0 U1816 ( .IN1(\regf[2][30] ), .IN2(n1401), .QN(n1769) );
  NAND2X0 U1817 ( .IN1(n1395), .IN2(\regf[1][0] ), .QN(n2355) );
  NAND2X0 U1818 ( .IN1(n1435), .IN2(\regf[1][0] ), .QN(n1888) );
  NAND2X0 U1819 ( .IN1(\regf[1][2] ), .IN2(n1389), .QN(n2347) );
  NAND2X0 U1820 ( .IN1(n1386), .IN2(\regf[1][3] ), .QN(n2343) );
  NAND2X0 U1821 ( .IN1(n1389), .IN2(\regf[1][31] ), .QN(n2231) );
  NAND2X0 U1822 ( .IN1(n1423), .IN2(\regf[1][2] ), .QN(n1880) );
  NAND2X0 U1823 ( .IN1(n1429), .IN2(\regf[1][3] ), .QN(n1876) );
  NAND2X0 U1824 ( .IN1(n1422), .IN2(\regf[1][31] ), .QN(n1764) );
  NAND2X0 U1825 ( .IN1(n1152), .IN2(\regf[1][1] ), .QN(n2351) );
  NAND2X0 U1826 ( .IN1(n1195), .IN2(\regf[1][1] ), .QN(n1884) );
  NAND2X0 U1827 ( .IN1(n1435), .IN2(\regf[1][20] ), .QN(n1808) );
  NAND2X0 U1828 ( .IN1(n1439), .IN2(\regf[1][21] ), .QN(n1804) );
  NAND2X0 U1829 ( .IN1(n1433), .IN2(\regf[1][22] ), .QN(n1800) );
  NAND2X0 U1830 ( .IN1(n1422), .IN2(\regf[1][23] ), .QN(n1796) );
  NAND2X0 U1831 ( .IN1(n1195), .IN2(\regf[1][24] ), .QN(n1792) );
  NAND2X0 U1832 ( .IN1(n1435), .IN2(\regf[1][25] ), .QN(n1788) );
  NAND2X0 U1833 ( .IN1(n1398), .IN2(\regf[1][26] ), .QN(n1784) );
  NAND2X0 U1834 ( .IN1(n1195), .IN2(\regf[1][27] ), .QN(n1780) );
  NAND2X0 U1835 ( .IN1(n1422), .IN2(\regf[1][28] ), .QN(n1776) );
  NAND2X0 U1836 ( .IN1(n1395), .IN2(\regf[1][5] ), .QN(n2335) );
  NAND2X0 U1837 ( .IN1(\regf[1][7] ), .IN2(n1103), .QN(n2327) );
  NAND2X0 U1838 ( .IN1(n1395), .IN2(\regf[1][8] ), .QN(n2323) );
  NAND2X0 U1839 ( .IN1(n1386), .IN2(\regf[1][9] ), .QN(n2319) );
  NAND2X0 U1840 ( .IN1(n1364), .IN2(\regf[1][10] ), .QN(n2315) );
  NAND2X0 U1841 ( .IN1(n1393), .IN2(\regf[1][11] ), .QN(n2311) );
  NAND2X0 U1842 ( .IN1(n1186), .IN2(\regf[1][12] ), .QN(n2307) );
  NAND2X0 U1843 ( .IN1(n1389), .IN2(\regf[1][13] ), .QN(n2303) );
  NAND2X0 U1844 ( .IN1(\regf[1][14] ), .IN2(n1371), .QN(n2299) );
  NAND2X0 U1845 ( .IN1(n1386), .IN2(\regf[1][15] ), .QN(n2295) );
  NAND2X0 U1846 ( .IN1(n1395), .IN2(\regf[1][16] ), .QN(n2291) );
  NAND2X0 U1847 ( .IN1(n1389), .IN2(\regf[1][17] ), .QN(n2287) );
  NAND2X0 U1848 ( .IN1(n1395), .IN2(\regf[1][18] ), .QN(n2283) );
  NAND2X0 U1849 ( .IN1(n1386), .IN2(\regf[1][19] ), .QN(n2279) );
  NAND2X0 U1850 ( .IN1(n1189), .IN2(\regf[1][20] ), .QN(n2275) );
  NAND2X0 U1851 ( .IN1(n1189), .IN2(\regf[1][21] ), .QN(n2271) );
  NAND2X0 U1852 ( .IN1(n1103), .IN2(\regf[1][22] ), .QN(n2267) );
  NAND2X0 U1853 ( .IN1(n1386), .IN2(\regf[1][23] ), .QN(n2263) );
  NAND2X0 U1854 ( .IN1(n1187), .IN2(\regf[1][24] ), .QN(n2259) );
  NAND2X0 U1855 ( .IN1(n1386), .IN2(\regf[1][25] ), .QN(n2255) );
  NAND2X0 U1856 ( .IN1(n1390), .IN2(\regf[1][26] ), .QN(n2251) );
  NAND2X0 U1857 ( .IN1(n1381), .IN2(\regf[1][27] ), .QN(n2247) );
  NAND2X0 U1858 ( .IN1(n1392), .IN2(\regf[1][28] ), .QN(n2243) );
  NAND2X0 U1859 ( .IN1(n1440), .IN2(\regf[1][5] ), .QN(n1868) );
  NAND2X0 U1860 ( .IN1(n1435), .IN2(\regf[1][7] ), .QN(n1860) );
  NAND2X0 U1861 ( .IN1(n1085), .IN2(\regf[1][8] ), .QN(n1856) );
  NAND2X0 U1862 ( .IN1(n1431), .IN2(\regf[1][9] ), .QN(n1852) );
  NAND2X0 U1863 ( .IN1(n1075), .IN2(\regf[1][10] ), .QN(n1848) );
  NAND2X0 U1864 ( .IN1(n1432), .IN2(\regf[1][11] ), .QN(n1844) );
  NAND2X0 U1865 ( .IN1(n1195), .IN2(\regf[1][12] ), .QN(n1840) );
  NAND2X0 U1866 ( .IN1(n1397), .IN2(\regf[1][13] ), .QN(n1836) );
  NAND2X0 U1867 ( .IN1(n1419), .IN2(\regf[1][14] ), .QN(n1832) );
  NAND2X0 U1868 ( .IN1(n1410), .IN2(\regf[1][15] ), .QN(n1828) );
  NAND2X0 U1869 ( .IN1(n1405), .IN2(\regf[1][16] ), .QN(n1824) );
  NAND2X0 U1870 ( .IN1(n1409), .IN2(\regf[1][17] ), .QN(n1820) );
  NAND2X0 U1871 ( .IN1(n1435), .IN2(\regf[1][18] ), .QN(n1816) );
  NAND2X0 U1872 ( .IN1(n1435), .IN2(\regf[1][19] ), .QN(n1812) );
  NAND2X0 U1873 ( .IN1(n1372), .IN2(\regf[1][4] ), .QN(n2339) );
  NAND2X0 U1874 ( .IN1(n1391), .IN2(\regf[1][6] ), .QN(n2331) );
  NAND2X0 U1875 ( .IN1(n1389), .IN2(\regf[1][29] ), .QN(n2239) );
  NAND2X0 U1876 ( .IN1(n1435), .IN2(\regf[1][4] ), .QN(n1872) );
  NAND2X0 U1877 ( .IN1(n1421), .IN2(\regf[1][6] ), .QN(n1864) );
  NAND2X0 U1878 ( .IN1(n1076), .IN2(\regf[1][29] ), .QN(n1772) );
  NAND2X0 U1879 ( .IN1(n1811), .IN2(n1810), .QN(n1652) );
  NAND2X0 U1880 ( .IN1(\regf[2][20] ), .IN2(n1406), .QN(n1809) );
  NAND2X0 U1881 ( .IN1(n1807), .IN2(n1806), .QN(n1662) );
  NAND2X0 U1882 ( .IN1(\regf[2][21] ), .IN2(n1406), .QN(n1805) );
  NAND2X0 U1883 ( .IN1(n1803), .IN2(n1802), .QN(n1672) );
  NAND2X0 U1884 ( .IN1(n1799), .IN2(n1798), .QN(n1682) );
  NAND2X0 U1885 ( .IN1(\regf[2][23] ), .IN2(n1403), .QN(n1797) );
  NAND2X0 U1886 ( .IN1(n1795), .IN2(n1794), .QN(n1692) );
  NAND2X0 U1887 ( .IN1(\regf[2][24] ), .IN2(n1399), .QN(n1793) );
  NAND2X0 U1888 ( .IN1(n1791), .IN2(n1790), .QN(n1702) );
  NAND2X0 U1889 ( .IN1(\regf[2][25] ), .IN2(n1406), .QN(n1789) );
  NAND2X0 U1890 ( .IN1(n1787), .IN2(n1786), .QN(n1712) );
  NAND2X0 U1891 ( .IN1(\regf[2][26] ), .IN2(n1408), .QN(n1785) );
  NAND2X0 U1892 ( .IN1(n1783), .IN2(n1782), .QN(n1722) );
  NAND2X0 U1893 ( .IN1(\regf[2][27] ), .IN2(n1401), .QN(n1781) );
  NAND2X0 U1894 ( .IN1(n1779), .IN2(n1778), .QN(n1732) );
  NAND2X0 U1895 ( .IN1(\regf[2][28] ), .IN2(n1408), .QN(n1777) );
  NAND2X0 U1896 ( .IN1(n2337), .IN2(n2338), .QN(n1969) );
  NAND2X0 U1897 ( .IN1(n2330), .IN2(n2329), .QN(n1989) );
  NAND2X0 U1898 ( .IN1(\regf[2][7] ), .IN2(n2363), .QN(n2328) );
  NAND2X0 U1899 ( .IN1(n2326), .IN2(n2325), .QN(n1999) );
  NAND2X0 U1900 ( .IN1(\regf[2][8] ), .IN2(n1360), .QN(n2324) );
  NAND2X0 U1901 ( .IN1(n2322), .IN2(n2321), .QN(n2009) );
  NAND2X0 U1902 ( .IN1(\regf[2][9] ), .IN2(n2363), .QN(n2320) );
  NAND2X0 U1903 ( .IN1(n2317), .IN2(n2318), .QN(n2019) );
  NAND2X0 U1904 ( .IN1(\regf[2][10] ), .IN2(n2365), .QN(n2316) );
  NAND2X0 U1905 ( .IN1(n2314), .IN2(n2313), .QN(n2029) );
  NAND2X0 U1906 ( .IN1(\regf[2][11] ), .IN2(n1360), .QN(n2312) );
  NAND2X0 U1907 ( .IN1(n2310), .IN2(n2309), .QN(n2039) );
  NAND2X0 U1908 ( .IN1(n2305), .IN2(n2306), .QN(n2049) );
  NAND2X0 U1909 ( .IN1(\regf[2][13] ), .IN2(n2365), .QN(n2304) );
  NAND2X0 U1910 ( .IN1(n2302), .IN2(n2301), .QN(n2059) );
  NAND2X0 U1911 ( .IN1(n2298), .IN2(n2297), .QN(n2069) );
  NAND2X0 U1912 ( .IN1(\regf[2][15] ), .IN2(n2364), .QN(n2296) );
  NAND2X0 U1913 ( .IN1(n2294), .IN2(n2293), .QN(n2079) );
  NAND2X0 U1914 ( .IN1(\regf[2][16] ), .IN2(n1361), .QN(n2292) );
  NAND2X0 U1915 ( .IN1(n2290), .IN2(n2289), .QN(n2089) );
  NAND2X0 U1916 ( .IN1(\regf[2][17] ), .IN2(n2363), .QN(n2288) );
  NAND2X0 U1917 ( .IN1(n2286), .IN2(n2285), .QN(n2099) );
  NAND2X0 U1918 ( .IN1(\regf[2][18] ), .IN2(n1361), .QN(n2284) );
  NAND2X0 U1919 ( .IN1(n2282), .IN2(n2281), .QN(n2109) );
  NAND2X0 U1920 ( .IN1(\regf[2][19] ), .IN2(n2363), .QN(n2280) );
  NAND2X0 U1921 ( .IN1(n2278), .IN2(n2277), .QN(n2119) );
  NAND2X0 U1922 ( .IN1(\regf[2][20] ), .IN2(n1361), .QN(n2276) );
  NAND2X0 U1923 ( .IN1(n2274), .IN2(n2273), .QN(n2129) );
  NAND2X0 U1924 ( .IN1(\regf[2][21] ), .IN2(n2363), .QN(n2272) );
  NAND2X0 U1925 ( .IN1(n2270), .IN2(n2269), .QN(n2139) );
  NAND2X0 U1926 ( .IN1(\regf[2][22] ), .IN2(n1361), .QN(n2268) );
  NAND2X0 U1927 ( .IN1(n2266), .IN2(n2265), .QN(n2149) );
  NAND2X0 U1928 ( .IN1(\regf[2][23] ), .IN2(n1361), .QN(n2264) );
  NAND2X0 U1929 ( .IN1(n2262), .IN2(n2261), .QN(n2159) );
  NAND2X0 U1930 ( .IN1(\regf[2][24] ), .IN2(n2362), .QN(n2260) );
  NAND2X0 U1931 ( .IN1(n2258), .IN2(n2257), .QN(n2169) );
  NAND2X0 U1932 ( .IN1(n2254), .IN2(n2253), .QN(n2179) );
  NAND2X0 U1933 ( .IN1(\regf[2][26] ), .IN2(n2365), .QN(n2252) );
  NAND2X0 U1934 ( .IN1(n2250), .IN2(n2249), .QN(n2189) );
  NAND2X0 U1935 ( .IN1(\regf[2][27] ), .IN2(n2364), .QN(n2248) );
  NAND2X0 U1936 ( .IN1(n2246), .IN2(n2245), .QN(n2199) );
  NAND2X0 U1937 ( .IN1(\regf[2][28] ), .IN2(n1360), .QN(n2244) );
  NAND2X0 U1938 ( .IN1(n1871), .IN2(n1870), .QN(n1502) );
  NAND2X0 U1939 ( .IN1(\regf[2][5] ), .IN2(n1401), .QN(n1869) );
  NAND2X0 U1940 ( .IN1(n1863), .IN2(n1862), .QN(n1522) );
  NAND2X0 U1941 ( .IN1(\regf[2][7] ), .IN2(n1893), .QN(n1861) );
  NAND2X0 U1942 ( .IN1(n1859), .IN2(n1858), .QN(n1532) );
  NAND2X0 U1943 ( .IN1(\regf[2][8] ), .IN2(n1893), .QN(n1857) );
  NAND2X0 U1944 ( .IN1(n1855), .IN2(n1854), .QN(n1542) );
  NAND2X0 U1945 ( .IN1(\regf[2][9] ), .IN2(n1399), .QN(n1853) );
  NAND2X0 U1946 ( .IN1(n1851), .IN2(n1850), .QN(n1552) );
  NAND2X0 U1947 ( .IN1(\regf[2][10] ), .IN2(n1893), .QN(n1849) );
  NAND2X0 U1948 ( .IN1(n1847), .IN2(n1846), .QN(n1562) );
  NAND2X0 U1949 ( .IN1(\regf[2][11] ), .IN2(n1408), .QN(n1845) );
  NAND2X0 U1950 ( .IN1(n1843), .IN2(n1842), .QN(n1572) );
  NAND2X0 U1951 ( .IN1(\regf[2][12] ), .IN2(n1399), .QN(n1841) );
  NAND2X0 U1952 ( .IN1(n1839), .IN2(n1838), .QN(n1582) );
  NAND2X0 U1953 ( .IN1(\regf[2][13] ), .IN2(n1406), .QN(n1837) );
  NAND2X0 U1954 ( .IN1(n1835), .IN2(n1834), .QN(n1592) );
  NAND2X0 U1955 ( .IN1(\regf[2][14] ), .IN2(n1893), .QN(n1833) );
  NAND2X0 U1956 ( .IN1(n1831), .IN2(n1830), .QN(n1602) );
  NAND2X0 U1957 ( .IN1(\regf[2][15] ), .IN2(n1893), .QN(n1829) );
  NAND2X0 U1958 ( .IN1(n1827), .IN2(n1826), .QN(n1612) );
  NAND2X0 U1959 ( .IN1(\regf[2][16] ), .IN2(n1406), .QN(n1825) );
  NAND2X0 U1960 ( .IN1(n1823), .IN2(n1822), .QN(n1622) );
  NAND2X0 U1961 ( .IN1(\regf[2][17] ), .IN2(n1408), .QN(n1821) );
  NAND2X0 U1962 ( .IN1(n1819), .IN2(n1818), .QN(n1632) );
  NAND2X0 U1963 ( .IN1(\regf[2][18] ), .IN2(n1893), .QN(n1817) );
  NAND2X0 U1964 ( .IN1(n1815), .IN2(n1814), .QN(n1642) );
  NAND2X0 U1965 ( .IN1(\regf[2][19] ), .IN2(n1401), .QN(n1813) );
  NAND2X0 U1966 ( .IN1(n2358), .IN2(n2357), .QN(n1919) );
  NAND2X0 U1967 ( .IN1(\regf[2][0] ), .IN2(n2364), .QN(n2356) );
  NAND2X0 U1968 ( .IN1(n1891), .IN2(n1890), .QN(n1452) );
  NAND2X0 U1969 ( .IN1(\regf[2][0] ), .IN2(n1406), .QN(n1889) );
  NAND2X0 U1970 ( .IN1(n2242), .IN2(n2241), .QN(n2209) );
  NAND2X0 U1971 ( .IN1(\regf[2][29] ), .IN2(n2366), .QN(n2240) );
  NAND2X0 U1972 ( .IN1(n1775), .IN2(n1774), .QN(n1742) );
  NAND2X0 U1973 ( .IN1(\regf[2][29] ), .IN2(n1399), .QN(n1773) );
  NAND2X0 U1974 ( .IN1(n2234), .IN2(n2233), .QN(n2229) );
  NAND2X0 U1975 ( .IN1(\regf[2][31] ), .IN2(n1360), .QN(n2232) );
  NAND2X0 U1976 ( .IN1(n1767), .IN2(n1766), .QN(n1762) );
  NAND2X0 U1977 ( .IN1(\regf[2][31] ), .IN2(n1893), .QN(n1765) );
  NAND2X0 U1978 ( .IN1(n2342), .IN2(n2341), .QN(n1959) );
  NAND2X0 U1979 ( .IN1(\regf[2][4] ), .IN2(n2364), .QN(n2340) );
  NAND2X0 U1980 ( .IN1(n2333), .IN2(n2334), .QN(n1979) );
  NAND2X0 U1981 ( .IN1(\regf[2][6] ), .IN2(n2365), .QN(n2332) );
  NAND2X0 U1982 ( .IN1(n1875), .IN2(n1874), .QN(n1492) );
  NAND2X0 U1983 ( .IN1(\regf[2][4] ), .IN2(n1408), .QN(n1873) );
  NAND2X0 U1984 ( .IN1(n1867), .IN2(n1866), .QN(n1512) );
  NAND2X0 U1985 ( .IN1(n2350), .IN2(n2349), .QN(n1939) );
  NAND2X0 U1986 ( .IN1(\regf[2][2] ), .IN2(n1360), .QN(n2348) );
  NAND2X0 U1987 ( .IN1(n2346), .IN2(n2345), .QN(n1949) );
  NAND2X0 U1988 ( .IN1(n1883), .IN2(n1882), .QN(n1472) );
  NAND2X0 U1989 ( .IN1(\regf[2][2] ), .IN2(n1401), .QN(n1881) );
  NAND2X0 U1990 ( .IN1(n1879), .IN2(n1878), .QN(n1482) );
  NAND2X0 U1991 ( .IN1(\regf[2][3] ), .IN2(n1406), .QN(n1877) );
  NAND2X0 U1992 ( .IN1(n2354), .IN2(n2353), .QN(n1929) );
  NAND2X0 U1993 ( .IN1(\regf[2][1] ), .IN2(n1361), .QN(n2352) );
  NAND2X0 U1994 ( .IN1(n1887), .IN2(n1886), .QN(n1462) );
  NBUFFX2 U1995 ( .INP(N19), .Z(n2374) );
  NBUFFX2 U1996 ( .INP(N14), .Z(n1902) );
  NBUFFX2 U1997 ( .INP(N20), .Z(n2381) );
  NBUFFX2 U1998 ( .INP(N15), .Z(n1909) );
  NBUFFX2 U1999 ( .INP(N19), .Z(n2375) );
  NBUFFX2 U2000 ( .INP(N19), .Z(n2376) );
  NBUFFX2 U2001 ( .INP(N19), .Z(n2377) );
  NBUFFX2 U2002 ( .INP(N19), .Z(n2378) );
  NBUFFX2 U2003 ( .INP(N14), .Z(n1903) );
  NBUFFX2 U2004 ( .INP(N14), .Z(n1904) );
  NBUFFX2 U2005 ( .INP(N14), .Z(n1905) );
  NBUFFX2 U2006 ( .INP(N20), .Z(n2380) );
  NBUFFX2 U2007 ( .INP(N15), .Z(n1908) );
  NBUFFX2 U2008 ( .INP(N18), .Z(n2368) );
  NBUFFX2 U2009 ( .INP(N13), .Z(n1896) );
  AND3X1 U2010 ( .IN1(wr_en), .IN2(n2711), .IN3(wr_addr[3]), .Q(n53) );
  INVX0 U2011 ( .INP(wr_addr[3]), .ZN(n2712) );
  NBUFFX2 U2012 ( .INP(wr_data[0]), .Z(n2525) );
  NBUFFX2 U2013 ( .INP(wr_data[1]), .Z(n2528) );
  NBUFFX2 U2014 ( .INP(wr_data[2]), .Z(n2531) );
  NBUFFX2 U2015 ( .INP(wr_data[3]), .Z(n2534) );
  NBUFFX2 U2016 ( .INP(wr_data[4]), .Z(n2537) );
  NBUFFX2 U2017 ( .INP(wr_data[5]), .Z(n2540) );
  NBUFFX2 U2018 ( .INP(wr_data[6]), .Z(n2543) );
  NBUFFX2 U2019 ( .INP(wr_data[7]), .Z(n2546) );
  NBUFFX2 U2020 ( .INP(wr_data[8]), .Z(n2549) );
  NBUFFX2 U2021 ( .INP(wr_data[9]), .Z(n2552) );
  NBUFFX2 U2022 ( .INP(wr_data[10]), .Z(n2555) );
  NBUFFX2 U2023 ( .INP(wr_data[11]), .Z(n2558) );
  NBUFFX2 U2024 ( .INP(wr_data[12]), .Z(n2561) );
  NBUFFX2 U2025 ( .INP(wr_data[13]), .Z(n2564) );
  NBUFFX2 U2026 ( .INP(wr_data[14]), .Z(n2567) );
  NBUFFX2 U2027 ( .INP(wr_data[15]), .Z(n2570) );
  NBUFFX2 U2028 ( .INP(wr_data[16]), .Z(n2573) );
  NBUFFX2 U2029 ( .INP(wr_data[17]), .Z(n2576) );
  NBUFFX2 U2030 ( .INP(wr_data[18]), .Z(n2579) );
  NBUFFX2 U2031 ( .INP(wr_data[19]), .Z(n2582) );
  NBUFFX2 U2032 ( .INP(wr_data[20]), .Z(n2585) );
  NBUFFX2 U2033 ( .INP(wr_data[21]), .Z(n2588) );
  NBUFFX2 U2034 ( .INP(wr_data[22]), .Z(n2591) );
  NBUFFX2 U2035 ( .INP(wr_data[23]), .Z(n2594) );
  NBUFFX2 U2036 ( .INP(wr_data[24]), .Z(n2597) );
  NBUFFX2 U2037 ( .INP(wr_data[25]), .Z(n2600) );
  NBUFFX2 U2038 ( .INP(wr_data[26]), .Z(n2603) );
  NBUFFX2 U2039 ( .INP(wr_data[27]), .Z(n2606) );
  NBUFFX2 U2040 ( .INP(wr_data[28]), .Z(n2609) );
  NBUFFX2 U2041 ( .INP(wr_data[29]), .Z(n2612) );
  NBUFFX2 U2042 ( .INP(wr_data[30]), .Z(n2615) );
  NBUFFX2 U2043 ( .INP(wr_data[31]), .Z(n2618) );
  NBUFFX2 U2044 ( .INP(wr_data[0]), .Z(n2526) );
  NBUFFX2 U2045 ( .INP(wr_data[1]), .Z(n2529) );
  NBUFFX2 U2046 ( .INP(wr_data[2]), .Z(n2532) );
  NBUFFX2 U2047 ( .INP(wr_data[3]), .Z(n2535) );
  NBUFFX2 U2048 ( .INP(wr_data[4]), .Z(n2538) );
  NBUFFX2 U2049 ( .INP(wr_data[5]), .Z(n2541) );
  NBUFFX2 U2050 ( .INP(wr_data[6]), .Z(n2544) );
  NBUFFX2 U2051 ( .INP(wr_data[7]), .Z(n2547) );
  NBUFFX2 U2052 ( .INP(wr_data[8]), .Z(n2550) );
  NBUFFX2 U2053 ( .INP(wr_data[9]), .Z(n2553) );
  NBUFFX2 U2054 ( .INP(wr_data[10]), .Z(n2556) );
  NBUFFX2 U2055 ( .INP(wr_data[11]), .Z(n2559) );
  NBUFFX2 U2056 ( .INP(wr_data[12]), .Z(n2562) );
  NBUFFX2 U2057 ( .INP(wr_data[13]), .Z(n2565) );
  NBUFFX2 U2058 ( .INP(wr_data[14]), .Z(n2568) );
  NBUFFX2 U2059 ( .INP(wr_data[15]), .Z(n2571) );
  NBUFFX2 U2060 ( .INP(wr_data[16]), .Z(n2574) );
  NBUFFX2 U2061 ( .INP(wr_data[17]), .Z(n2577) );
  NBUFFX2 U2062 ( .INP(wr_data[18]), .Z(n2580) );
  NBUFFX2 U2063 ( .INP(wr_data[19]), .Z(n2583) );
  NBUFFX2 U2064 ( .INP(wr_data[20]), .Z(n2586) );
  NBUFFX2 U2065 ( .INP(wr_data[21]), .Z(n2589) );
  NBUFFX2 U2066 ( .INP(wr_data[22]), .Z(n2592) );
  NBUFFX2 U2067 ( .INP(wr_data[23]), .Z(n2595) );
  NBUFFX2 U2068 ( .INP(wr_data[24]), .Z(n2598) );
  NBUFFX2 U2069 ( .INP(wr_data[25]), .Z(n2601) );
  NBUFFX2 U2070 ( .INP(wr_data[26]), .Z(n2604) );
  NBUFFX2 U2071 ( .INP(wr_data[27]), .Z(n2607) );
  NBUFFX2 U2072 ( .INP(wr_data[28]), .Z(n2610) );
  NBUFFX2 U2073 ( .INP(wr_data[29]), .Z(n2613) );
  NBUFFX2 U2074 ( .INP(wr_data[30]), .Z(n2616) );
  NBUFFX2 U2075 ( .INP(wr_data[31]), .Z(n2619) );
  NBUFFX2 U2076 ( .INP(wr_data[0]), .Z(n2527) );
  NBUFFX2 U2077 ( .INP(wr_data[1]), .Z(n2530) );
  NBUFFX2 U2078 ( .INP(wr_data[2]), .Z(n2533) );
  NBUFFX2 U2079 ( .INP(wr_data[3]), .Z(n2536) );
  NBUFFX2 U2080 ( .INP(wr_data[14]), .Z(n2569) );
  NBUFFX2 U2081 ( .INP(wr_data[15]), .Z(n2572) );
  NBUFFX2 U2082 ( .INP(wr_data[16]), .Z(n2575) );
  NBUFFX2 U2083 ( .INP(wr_data[17]), .Z(n2578) );
  NBUFFX2 U2084 ( .INP(wr_data[18]), .Z(n2581) );
  NBUFFX2 U2085 ( .INP(wr_data[19]), .Z(n2584) );
  NBUFFX2 U2086 ( .INP(wr_data[4]), .Z(n2539) );
  NBUFFX2 U2087 ( .INP(wr_data[5]), .Z(n2542) );
  NBUFFX2 U2088 ( .INP(wr_data[6]), .Z(n2545) );
  NBUFFX2 U2089 ( .INP(wr_data[7]), .Z(n2548) );
  NBUFFX2 U2090 ( .INP(wr_data[8]), .Z(n2551) );
  NBUFFX2 U2091 ( .INP(wr_data[9]), .Z(n2554) );
  NBUFFX2 U2092 ( .INP(wr_data[10]), .Z(n2557) );
  NBUFFX2 U2093 ( .INP(wr_data[11]), .Z(n2560) );
  NBUFFX2 U2094 ( .INP(wr_data[12]), .Z(n2563) );
  NBUFFX2 U2095 ( .INP(wr_data[13]), .Z(n2566) );
  NBUFFX2 U2096 ( .INP(wr_data[20]), .Z(n2587) );
  NBUFFX2 U2097 ( .INP(wr_data[21]), .Z(n2590) );
  NBUFFX2 U2098 ( .INP(wr_data[22]), .Z(n2593) );
  NBUFFX2 U2099 ( .INP(wr_data[23]), .Z(n2596) );
  NBUFFX2 U2100 ( .INP(wr_data[24]), .Z(n2599) );
  NBUFFX2 U2101 ( .INP(wr_data[25]), .Z(n2602) );
  NBUFFX2 U2102 ( .INP(wr_data[26]), .Z(n2605) );
  NBUFFX2 U2103 ( .INP(wr_data[27]), .Z(n2608) );
  NBUFFX2 U2104 ( .INP(wr_data[28]), .Z(n2611) );
  NBUFFX2 U2105 ( .INP(wr_data[29]), .Z(n2614) );
  NBUFFX2 U2106 ( .INP(wr_data[30]), .Z(n2617) );
  NBUFFX2 U2107 ( .INP(wr_data[31]), .Z(n2620) );
  NBUFFX2 U2108 ( .INP(nrst), .Z(n2704) );
  NBUFFX2 U2109 ( .INP(nrst), .Z(n2705) );
  NBUFFX2 U2110 ( .INP(nrst), .Z(n2706) );
  NBUFFX2 U2111 ( .INP(nrst), .Z(n2707) );
  NBUFFX2 U2112 ( .INP(nrst), .Z(n2708) );
  NBUFFX2 U2113 ( .INP(nrst), .Z(n2709) );
  NBUFFX2 U2114 ( .INP(nrst), .Z(n2710) );
  MUX41X1 U2115 ( .IN1(\regf[28][0] ), .IN3(\regf[30][0] ), .IN2(\regf[29][0] ), .IN4(\regf[31][0] ), .S0(n1287), .S1(n1197), .Q(n1444) );
  MUX41X1 U2116 ( .IN1(\regf[24][0] ), .IN3(\regf[26][0] ), .IN2(\regf[25][0] ), .IN4(\regf[27][0] ), .S0(n1348), .S1(n1185), .Q(n1445) );
  MUX41X1 U2117 ( .IN1(\regf[16][0] ), .IN3(\regf[18][0] ), .IN2(\regf[17][0] ), .IN4(\regf[19][0] ), .S0(n1344), .S1(n1428), .Q(n1447) );
  MUX41X1 U2118 ( .IN1(n1447), .IN3(n1445), .IN2(n1446), .IN4(n1444), .S0(
        n1902), .S1(n1896), .Q(n1448) );
  MUX41X1 U2119 ( .IN1(\regf[12][0] ), .IN3(\regf[14][0] ), .IN2(\regf[13][0] ), .IN4(\regf[15][0] ), .S0(n1349), .S1(n1440), .Q(n1449) );
  MUX41X1 U2120 ( .IN1(\regf[8][0] ), .IN3(\regf[10][0] ), .IN2(\regf[9][0] ), 
        .IN4(\regf[11][0] ), .S0(n1293), .S1(n1119), .Q(n1450) );
  MUX41X1 U2121 ( .IN1(\regf[4][0] ), .IN3(\regf[6][0] ), .IN2(\regf[5][0] ), 
        .IN4(\regf[7][0] ), .S0(n1344), .S1(n1158), .Q(n1451) );
  MUX41X1 U2122 ( .IN1(n1452), .IN3(n1450), .IN2(n1451), .IN4(n1449), .S0(
        n1902), .S1(n1896), .Q(n1453) );
  MUX41X1 U2123 ( .IN1(\regf[28][1] ), .IN3(\regf[30][1] ), .IN2(\regf[29][1] ), .IN4(\regf[31][1] ), .S0(n1345), .S1(n1397), .Q(n1454) );
  MUX41X1 U2124 ( .IN1(\regf[24][1] ), .IN3(\regf[26][1] ), .IN2(\regf[25][1] ), .IN4(\regf[27][1] ), .S0(n1285), .S1(n1418), .Q(n1455) );
  MUX41X1 U2125 ( .IN1(\regf[20][1] ), .IN3(\regf[22][1] ), .IN2(\regf[21][1] ), .IN4(\regf[23][1] ), .S0(n1349), .S1(n1428), .Q(n1456) );
  MUX41X1 U2126 ( .IN1(\regf[16][1] ), .IN3(\regf[18][1] ), .IN2(\regf[17][1] ), .IN4(\regf[19][1] ), .S0(n1285), .S1(n1421), .Q(n1457) );
  MUX41X1 U2127 ( .IN1(n1457), .IN3(n1455), .IN2(n1456), .IN4(n1454), .S0(
        n1902), .S1(n1896), .Q(n1458) );
  MUX41X1 U2128 ( .IN1(\regf[12][1] ), .IN3(\regf[14][1] ), .IN2(\regf[13][1] ), .IN4(\regf[15][1] ), .S0(n1350), .S1(n1428), .Q(n1459) );
  MUX41X1 U2129 ( .IN1(\regf[8][1] ), .IN3(\regf[10][1] ), .IN2(\regf[9][1] ), 
        .IN4(\regf[11][1] ), .S0(n1294), .S1(n1084), .Q(n1460) );
  MUX41X1 U2130 ( .IN1(\regf[4][1] ), .IN3(\regf[6][1] ), .IN2(\regf[5][1] ), 
        .IN4(\regf[7][1] ), .S0(n1345), .S1(n1180), .Q(n1461) );
  MUX21X1 U2131 ( .IN1(n1463), .IN2(n1458), .S(n1908), .Q(rd_dataA[1]) );
  MUX41X1 U2132 ( .IN1(\regf[28][2] ), .IN3(\regf[30][2] ), .IN2(\regf[29][2] ), .IN4(\regf[31][2] ), .S0(n1284), .S1(n1146), .Q(n1464) );
  MUX41X1 U2133 ( .IN1(\regf[24][2] ), .IN3(\regf[26][2] ), .IN2(\regf[25][2] ), .IN4(\regf[27][2] ), .S0(n1286), .S1(n1101), .Q(n1465) );
  MUX41X1 U2134 ( .IN1(\regf[20][2] ), .IN3(\regf[22][2] ), .IN2(\regf[21][2] ), .IN4(\regf[23][2] ), .S0(n1350), .S1(n1434), .Q(n1466) );
  MUX41X1 U2135 ( .IN1(\regf[16][2] ), .IN3(\regf[18][2] ), .IN2(\regf[17][2] ), .IN4(\regf[19][2] ), .S0(n1346), .S1(n1149), .Q(n1467) );
  MUX41X1 U2136 ( .IN1(n1467), .IN3(n1465), .IN2(n1466), .IN4(n1464), .S0(
        n1903), .S1(n1897), .Q(n1468) );
  MUX41X1 U2137 ( .IN1(\regf[8][2] ), .IN3(\regf[10][2] ), .IN2(\regf[9][2] ), 
        .IN4(\regf[11][2] ), .S0(n1317), .S1(n1114), .Q(n1470) );
  MUX41X1 U2138 ( .IN1(\regf[4][2] ), .IN3(\regf[6][2] ), .IN2(\regf[5][2] ), 
        .IN4(\regf[7][2] ), .S0(n1299), .S1(n1150), .Q(n1471) );
  MUX41X1 U2139 ( .IN1(n1472), .IN3(n1470), .IN2(n1471), .IN4(n1469), .S0(
        n1903), .S1(n1897), .Q(n1473) );
  MUX21X1 U2140 ( .IN1(n1473), .IN2(n1468), .S(n1908), .Q(rd_dataA[2]) );
  MUX41X1 U2141 ( .IN1(\regf[28][3] ), .IN3(\regf[30][3] ), .IN2(\regf[29][3] ), .IN4(\regf[31][3] ), .S0(n1334), .S1(n1402), .Q(n1474) );
  MUX41X1 U2142 ( .IN1(\regf[24][3] ), .IN3(\regf[26][3] ), .IN2(\regf[25][3] ), .IN4(\regf[27][3] ), .S0(n1288), .S1(n1443), .Q(n1475) );
  MUX41X1 U2143 ( .IN1(\regf[20][3] ), .IN3(\regf[22][3] ), .IN2(\regf[21][3] ), .IN4(\regf[23][3] ), .S0(n1337), .S1(n1410), .Q(n1476) );
  MUX41X1 U2144 ( .IN1(\regf[16][3] ), .IN3(\regf[18][3] ), .IN2(\regf[17][3] ), .IN4(\regf[19][3] ), .S0(n1134), .S1(n1146), .Q(n1477) );
  MUX41X1 U2145 ( .IN1(n1477), .IN3(n1475), .IN2(n1476), .IN4(n1474), .S0(
        n1903), .S1(n1897), .Q(n1478) );
  MUX41X1 U2146 ( .IN1(\regf[12][3] ), .IN3(\regf[14][3] ), .IN2(\regf[13][3] ), .IN4(\regf[15][3] ), .S0(n1290), .S1(n1074), .Q(n1479) );
  MUX41X1 U2147 ( .IN1(\regf[8][3] ), .IN3(\regf[10][3] ), .IN2(\regf[9][3] ), 
        .IN4(\regf[11][3] ), .S0(n1318), .S1(n1159), .Q(n1480) );
  MUX41X1 U2148 ( .IN1(\regf[4][3] ), .IN3(\regf[6][3] ), .IN2(\regf[5][3] ), 
        .IN4(\regf[7][3] ), .S0(n1300), .S1(n1437), .Q(n1481) );
  MUX21X1 U2149 ( .IN1(n1483), .IN2(n1478), .S(n1908), .Q(rd_dataA[3]) );
  MUX41X1 U2150 ( .IN1(\regf[28][4] ), .IN3(\regf[30][4] ), .IN2(\regf[29][4] ), .IN4(\regf[31][4] ), .S0(n1336), .S1(n1081), .Q(n1484) );
  MUX41X1 U2151 ( .IN1(\regf[24][4] ), .IN3(\regf[26][4] ), .IN2(\regf[25][4] ), .IN4(\regf[27][4] ), .S0(n1341), .S1(n1084), .Q(n1485) );
  MUX41X1 U2152 ( .IN1(\regf[20][4] ), .IN3(\regf[22][4] ), .IN2(\regf[21][4] ), .IN4(\regf[23][4] ), .S0(n1338), .S1(n1404), .Q(n1486) );
  MUX41X1 U2153 ( .IN1(\regf[16][4] ), .IN3(\regf[18][4] ), .IN2(\regf[17][4] ), .IN4(\regf[19][4] ), .S0(n1333), .S1(n1146), .Q(n1487) );
  MUX41X1 U2154 ( .IN1(n1487), .IN3(n1485), .IN2(n1486), .IN4(n1484), .S0(
        n1903), .S1(n1897), .Q(n1488) );
  MUX41X1 U2155 ( .IN1(\regf[12][4] ), .IN3(\regf[14][4] ), .IN2(\regf[13][4] ), .IN4(\regf[15][4] ), .S0(n1341), .S1(n1173), .Q(n1489) );
  MUX41X1 U2156 ( .IN1(\regf[8][4] ), .IN3(\regf[10][4] ), .IN2(\regf[9][4] ), 
        .IN4(\regf[11][4] ), .S0(n1319), .S1(n1150), .Q(n1490) );
  MUX41X1 U2157 ( .IN1(\regf[4][4] ), .IN3(\regf[6][4] ), .IN2(\regf[5][4] ), 
        .IN4(\regf[7][4] ), .S0(n1290), .S1(n1410), .Q(n1491) );
  MUX41X1 U2158 ( .IN1(n1492), .IN3(n1490), .IN2(n1491), .IN4(n1489), .S0(
        n1903), .S1(n1897), .Q(n1493) );
  MUX21X1 U2159 ( .IN1(n1493), .IN2(n1488), .S(n1908), .Q(rd_dataA[4]) );
  MUX41X1 U2160 ( .IN1(\regf[24][5] ), .IN3(\regf[26][5] ), .IN2(\regf[25][5] ), .IN4(\regf[27][5] ), .S0(n1288), .S1(n1073), .Q(n1495) );
  MUX41X1 U2161 ( .IN1(\regf[20][5] ), .IN3(\regf[22][5] ), .IN2(\regf[21][5] ), .IN4(\regf[23][5] ), .S0(n1290), .S1(n1431), .Q(n1496) );
  MUX41X1 U2162 ( .IN1(\regf[16][5] ), .IN3(\regf[18][5] ), .IN2(\regf[17][5] ), .IN4(\regf[19][5] ), .S0(n1329), .S1(n1423), .Q(n1497) );
  MUX41X1 U2163 ( .IN1(n1497), .IN3(n1495), .IN2(n1496), .IN4(n1494), .S0(
        n1903), .S1(n1897), .Q(n1498) );
  MUX41X1 U2164 ( .IN1(\regf[12][5] ), .IN3(\regf[14][5] ), .IN2(\regf[13][5] ), .IN4(\regf[15][5] ), .S0(n1283), .S1(n1433), .Q(n1499) );
  MUX41X1 U2165 ( .IN1(\regf[8][5] ), .IN3(\regf[10][5] ), .IN2(\regf[9][5] ), 
        .IN4(\regf[11][5] ), .S0(n1307), .S1(n1431), .Q(n1500) );
  MUX41X1 U2166 ( .IN1(\regf[4][5] ), .IN3(\regf[6][5] ), .IN2(\regf[5][5] ), 
        .IN4(\regf[7][5] ), .S0(n1304), .S1(n1405), .Q(n1501) );
  MUX41X1 U2167 ( .IN1(n1502), .IN3(n1500), .IN2(n1501), .IN4(n1499), .S0(
        n1903), .S1(n1897), .Q(n1503) );
  MUX41X1 U2168 ( .IN1(\regf[28][6] ), .IN3(\regf[30][6] ), .IN2(\regf[29][6] ), .IN4(\regf[31][6] ), .S0(n1288), .S1(n1419), .Q(n1504) );
  MUX41X1 U2169 ( .IN1(\regf[24][6] ), .IN3(\regf[26][6] ), .IN2(\regf[25][6] ), .IN4(\regf[27][6] ), .S0(n1339), .S1(n1427), .Q(n1505) );
  MUX41X1 U2170 ( .IN1(\regf[20][6] ), .IN3(\regf[22][6] ), .IN2(\regf[21][6] ), .IN4(\regf[23][6] ), .S0(n1346), .S1(n1146), .Q(n1506) );
  MUX41X1 U2171 ( .IN1(\regf[16][6] ), .IN3(\regf[18][6] ), .IN2(\regf[17][6] ), .IN4(\regf[19][6] ), .S0(n1330), .S1(n1432), .Q(n1507) );
  MUX41X1 U2172 ( .IN1(n1507), .IN3(n1505), .IN2(n1506), .IN4(n1504), .S0(
        n1903), .S1(n1897), .Q(n1508) );
  MUX41X1 U2173 ( .IN1(\regf[12][6] ), .IN3(\regf[14][6] ), .IN2(\regf[13][6] ), .IN4(\regf[15][6] ), .S0(n1339), .S1(n1082), .Q(n1509) );
  MUX41X1 U2174 ( .IN1(\regf[8][6] ), .IN3(\regf[10][6] ), .IN2(\regf[9][6] ), 
        .IN4(\regf[11][6] ), .S0(n1308), .S1(n1421), .Q(n1510) );
  MUX41X1 U2175 ( .IN1(\regf[4][6] ), .IN3(\regf[6][6] ), .IN2(\regf[5][6] ), 
        .IN4(\regf[7][6] ), .S0(n1305), .S1(n1176), .Q(n1511) );
  MUX41X1 U2176 ( .IN1(\regf[28][7] ), .IN3(\regf[30][7] ), .IN2(\regf[29][7] ), .IN4(\regf[31][7] ), .S0(n1319), .S1(n1441), .Q(n1514) );
  MUX41X1 U2177 ( .IN1(\regf[24][7] ), .IN3(\regf[26][7] ), .IN2(\regf[25][7] ), .IN4(\regf[27][7] ), .S0(n1338), .S1(n1423), .Q(n1515) );
  MUX41X1 U2178 ( .IN1(\regf[20][7] ), .IN3(\regf[22][7] ), .IN2(\regf[21][7] ), .IN4(\regf[23][7] ), .S0(n1344), .S1(n1397), .Q(n1516) );
  MUX41X1 U2179 ( .IN1(\regf[16][7] ), .IN3(\regf[18][7] ), .IN2(\regf[17][7] ), .IN4(\regf[19][7] ), .S0(n1325), .S1(n1405), .Q(n1517) );
  MUX41X1 U2180 ( .IN1(n1517), .IN3(n1515), .IN2(n1516), .IN4(n1514), .S0(
        n1903), .S1(n1897), .Q(n1518) );
  MUX41X1 U2181 ( .IN1(\regf[12][7] ), .IN3(\regf[14][7] ), .IN2(\regf[13][7] ), .IN4(\regf[15][7] ), .S0(n1337), .S1(n1430), .Q(n1519) );
  MUX41X1 U2182 ( .IN1(\regf[8][7] ), .IN3(\regf[10][7] ), .IN2(\regf[9][7] ), 
        .IN4(\regf[11][7] ), .S0(n1305), .S1(n1132), .Q(n1520) );
  MUX41X1 U2183 ( .IN1(\regf[4][7] ), .IN3(\regf[6][7] ), .IN2(\regf[5][7] ), 
        .IN4(\regf[7][7] ), .S0(n1288), .S1(n1079), .Q(n1521) );
  MUX41X1 U2184 ( .IN1(n1522), .IN3(n1520), .IN2(n1521), .IN4(n1519), .S0(
        n1903), .S1(n1897), .Q(n1523) );
  MUX21X1 U2185 ( .IN1(n1523), .IN2(n1518), .S(n1908), .Q(rd_dataA[7]) );
  MUX41X1 U2186 ( .IN1(\regf[28][8] ), .IN3(\regf[30][8] ), .IN2(\regf[29][8] ), .IN4(\regf[31][8] ), .S0(n1326), .S1(n1192), .Q(n1524) );
  MUX41X1 U2187 ( .IN1(\regf[24][8] ), .IN3(\regf[26][8] ), .IN2(\regf[25][8] ), .IN4(\regf[27][8] ), .S0(n1287), .S1(n1433), .Q(n1525) );
  MUX41X1 U2188 ( .IN1(\regf[20][8] ), .IN3(\regf[22][8] ), .IN2(\regf[21][8] ), .IN4(\regf[23][8] ), .S0(n1345), .S1(n1076), .Q(n1526) );
  MUX41X1 U2189 ( .IN1(\regf[16][8] ), .IN3(\regf[18][8] ), .IN2(\regf[17][8] ), .IN4(\regf[19][8] ), .S0(n1286), .S1(n1439), .Q(n1527) );
  MUX41X1 U2190 ( .IN1(n1527), .IN3(n1525), .IN2(n1526), .IN4(n1524), .S0(
        n1904), .S1(n1898), .Q(n1528) );
  MUX41X1 U2191 ( .IN1(\regf[12][8] ), .IN3(\regf[14][8] ), .IN2(\regf[13][8] ), .IN4(\regf[15][8] ), .S0(n1338), .S1(n1429), .Q(n1529) );
  MUX41X1 U2192 ( .IN1(\regf[8][8] ), .IN3(\regf[10][8] ), .IN2(\regf[9][8] ), 
        .IN4(\regf[11][8] ), .S0(n1306), .S1(n1178), .Q(n1530) );
  MUX41X1 U2193 ( .IN1(\regf[4][8] ), .IN3(\regf[6][8] ), .IN2(\regf[5][8] ), 
        .IN4(\regf[7][8] ), .S0(n1289), .S1(n1128), .Q(n1531) );
  MUX41X1 U2194 ( .IN1(n1532), .IN3(n1530), .IN2(n1531), .IN4(n1529), .S0(
        n1904), .S1(n1898), .Q(n1533) );
  MUX21X1 U2195 ( .IN1(n1533), .IN2(n1528), .S(n1909), .Q(rd_dataA[8]) );
  MUX41X1 U2196 ( .IN1(\regf[28][9] ), .IN3(\regf[30][9] ), .IN2(\regf[29][9] ), .IN4(\regf[31][9] ), .S0(n1327), .S1(n1427), .Q(n1534) );
  MUX41X1 U2197 ( .IN1(\regf[24][9] ), .IN3(\regf[26][9] ), .IN2(\regf[25][9] ), .IN4(\regf[27][9] ), .S0(n1331), .S1(n1183), .Q(n1535) );
  MUX41X1 U2198 ( .IN1(\regf[20][9] ), .IN3(\regf[22][9] ), .IN2(\regf[21][9] ), .IN4(\regf[23][9] ), .S0(n1285), .S1(n1430), .Q(n1536) );
  MUX41X1 U2199 ( .IN1(\regf[16][9] ), .IN3(\regf[18][9] ), .IN2(\regf[17][9] ), .IN4(\regf[19][9] ), .S0(n1307), .S1(n1075), .Q(n1537) );
  MUX41X1 U2200 ( .IN1(\regf[12][9] ), .IN3(\regf[14][9] ), .IN2(\regf[13][9] ), .IN4(\regf[15][9] ), .S0(n1331), .S1(n1085), .Q(n1539) );
  MUX41X1 U2201 ( .IN1(\regf[8][9] ), .IN3(\regf[10][9] ), .IN2(\regf[9][9] ), 
        .IN4(\regf[11][9] ), .S0(n1297), .S1(n1101), .Q(n1540) );
  MUX41X1 U2202 ( .IN1(\regf[4][9] ), .IN3(\regf[6][9] ), .IN2(\regf[5][9] ), 
        .IN4(\regf[7][9] ), .S0(n1288), .S1(n1129), .Q(n1541) );
  MUX41X1 U2203 ( .IN1(n1542), .IN3(n1540), .IN2(n1541), .IN4(n1539), .S0(
        n1904), .S1(n1898), .Q(n1543) );
  MUX21X1 U2204 ( .IN1(n1543), .IN2(n1538), .S(n1909), .Q(rd_dataA[9]) );
  MUX41X1 U2205 ( .IN1(\regf[28][10] ), .IN3(\regf[30][10] ), .IN2(
        \regf[29][10] ), .IN4(\regf[31][10] ), .S0(n1308), .S1(n1443), .Q(
        n1544) );
  MUX41X1 U2206 ( .IN1(\regf[24][10] ), .IN3(\regf[26][10] ), .IN2(
        \regf[25][10] ), .IN4(\regf[27][10] ), .S0(n1334), .S1(n1177), .Q(
        n1545) );
  MUX41X1 U2207 ( .IN1(\regf[20][10] ), .IN3(\regf[22][10] ), .IN2(
        \regf[21][10] ), .IN4(\regf[23][10] ), .S0(n1339), .S1(n1075), .Q(
        n1546) );
  MUX41X1 U2208 ( .IN1(\regf[16][10] ), .IN3(\regf[18][10] ), .IN2(
        \regf[17][10] ), .IN4(\regf[19][10] ), .S0(n1309), .S1(n1430), .Q(
        n1547) );
  MUX41X1 U2209 ( .IN1(n1547), .IN3(n1545), .IN2(n1546), .IN4(n1544), .S0(
        n1904), .S1(n1898), .Q(n1548) );
  MUX41X1 U2210 ( .IN1(\regf[12][10] ), .IN3(\regf[14][10] ), .IN2(
        \regf[13][10] ), .IN4(\regf[15][10] ), .S0(n1332), .S1(n1084), .Q(
        n1549) );
  MUX41X1 U2211 ( .IN1(\regf[8][10] ), .IN3(\regf[10][10] ), .IN2(
        \regf[9][10] ), .IN4(\regf[11][10] ), .S0(n1298), .S1(n1085), .Q(n1550) );
  MUX41X1 U2212 ( .IN1(\regf[4][10] ), .IN3(\regf[6][10] ), .IN2(\regf[5][10] ), .IN4(\regf[7][10] ), .S0(n1283), .S1(n1121), .Q(n1551) );
  MUX41X1 U2213 ( .IN1(n1552), .IN3(n1550), .IN2(n1551), .IN4(n1549), .S0(
        n1904), .S1(n1898), .Q(n1553) );
  MUX41X1 U2214 ( .IN1(\regf[28][11] ), .IN3(\regf[30][11] ), .IN2(
        \regf[29][11] ), .IN4(\regf[31][11] ), .S0(n1330), .S1(n1436), .Q(
        n1554) );
  MUX41X1 U2215 ( .IN1(\regf[24][11] ), .IN3(\regf[26][11] ), .IN2(
        \regf[25][11] ), .IN4(\regf[27][11] ), .S0(n1336), .S1(n1176), .Q(
        n1555) );
  MUX41X1 U2216 ( .IN1(\regf[16][11] ), .IN3(\regf[18][11] ), .IN2(
        \regf[17][11] ), .IN4(\regf[19][11] ), .S0(n1316), .S1(n1434), .Q(
        n1557) );
  MUX41X1 U2217 ( .IN1(n1557), .IN3(n1555), .IN2(n1556), .IN4(n1554), .S0(
        n1904), .S1(n1898), .Q(n1558) );
  MUX41X1 U2218 ( .IN1(\regf[12][11] ), .IN3(\regf[14][11] ), .IN2(
        \regf[13][11] ), .IN4(\regf[15][11] ), .S0(n1333), .S1(n1082), .Q(
        n1559) );
  MUX41X1 U2219 ( .IN1(\regf[8][11] ), .IN3(\regf[10][11] ), .IN2(
        \regf[9][11] ), .IN4(\regf[11][11] ), .S0(n1303), .S1(n1085), .Q(n1560) );
  MUX41X1 U2220 ( .IN1(\regf[4][11] ), .IN3(\regf[6][11] ), .IN2(\regf[5][11] ), .IN4(\regf[7][11] ), .S0(n1286), .S1(n1119), .Q(n1561) );
  MUX41X1 U2221 ( .IN1(n1562), .IN3(n1560), .IN2(n1561), .IN4(n1559), .S0(
        n1904), .S1(n1898), .Q(n1563) );
  MUX41X1 U2222 ( .IN1(\regf[28][12] ), .IN3(\regf[30][12] ), .IN2(
        \regf[29][12] ), .IN4(\regf[31][12] ), .S0(n1317), .S1(n1434), .Q(
        n1564) );
  MUX41X1 U2223 ( .IN1(\regf[20][12] ), .IN3(\regf[22][12] ), .IN2(
        \regf[21][12] ), .IN4(\regf[23][12] ), .S0(n1343), .S1(n1432), .Q(
        n1566) );
  MUX41X1 U2224 ( .IN1(n1567), .IN3(n1565), .IN2(n1566), .IN4(n1564), .S0(
        n1904), .S1(n1898), .Q(n1568) );
  MUX41X1 U2225 ( .IN1(\regf[12][12] ), .IN3(\regf[14][12] ), .IN2(
        \regf[13][12] ), .IN4(\regf[15][12] ), .S0(n1336), .S1(n1111), .Q(
        n1569) );
  MUX41X1 U2226 ( .IN1(\regf[8][12] ), .IN3(\regf[10][12] ), .IN2(
        \regf[9][12] ), .IN4(\regf[11][12] ), .S0(n1304), .S1(n1438), .Q(n1570) );
  MUX41X1 U2227 ( .IN1(\regf[4][12] ), .IN3(\regf[6][12] ), .IN2(\regf[5][12] ), .IN4(\regf[7][12] ), .S0(n1287), .S1(n1161), .Q(n1571) );
  MUX41X1 U2228 ( .IN1(n1572), .IN3(n1570), .IN2(n1571), .IN4(n1569), .S0(
        n1904), .S1(n1898), .Q(n1573) );
  MUX41X1 U2229 ( .IN1(\regf[28][13] ), .IN3(\regf[30][13] ), .IN2(
        \regf[29][13] ), .IN4(\regf[31][13] ), .S0(n1318), .S1(n1410), .Q(
        n1574) );
  MUX41X1 U2230 ( .IN1(\regf[24][13] ), .IN3(\regf[26][13] ), .IN2(
        \regf[25][13] ), .IN4(\regf[27][13] ), .S0(n1337), .S1(n1124), .Q(
        n1575) );
  MUX41X1 U2231 ( .IN1(\regf[20][13] ), .IN3(\regf[22][13] ), .IN2(
        \regf[21][13] ), .IN4(\regf[23][13] ), .S0(n1348), .S1(n1432), .Q(
        n1576) );
  MUX41X1 U2232 ( .IN1(\regf[12][13] ), .IN3(\regf[14][13] ), .IN2(
        \regf[13][13] ), .IN4(\regf[15][13] ), .S0(n1334), .S1(n1409), .Q(
        n1579) );
  MUX41X1 U2233 ( .IN1(\regf[8][13] ), .IN3(\regf[10][13] ), .IN2(
        \regf[9][13] ), .IN4(\regf[11][13] ), .S0(n1300), .S1(n1405), .Q(n1580) );
  MUX41X1 U2234 ( .IN1(\regf[4][13] ), .IN3(\regf[6][13] ), .IN2(\regf[5][13] ), .IN4(\regf[7][13] ), .S0(n1284), .S1(n1159), .Q(n1581) );
  MUX41X1 U2235 ( .IN1(n1582), .IN3(n1580), .IN2(n1581), .IN4(n1579), .S0(
        n1904), .S1(n1898), .Q(n1583) );
  MUX41X1 U2236 ( .IN1(\regf[28][14] ), .IN3(\regf[30][14] ), .IN2(
        \regf[29][14] ), .IN4(\regf[31][14] ), .S0(n1314), .S1(n1160), .Q(
        n1584) );
  MUX41X1 U2237 ( .IN1(\regf[20][14] ), .IN3(\regf[22][14] ), .IN2(
        \regf[21][14] ), .IN4(\regf[23][14] ), .S0(n1286), .S1(n1430), .Q(
        n1586) );
  MUX41X1 U2238 ( .IN1(\regf[16][14] ), .IN3(\regf[18][14] ), .IN2(
        \regf[17][14] ), .IN4(\regf[19][14] ), .S0(n1315), .S1(n1429), .Q(
        n1587) );
  MUX41X1 U2239 ( .IN1(\regf[12][14] ), .IN3(\regf[14][14] ), .IN2(
        \regf[13][14] ), .IN4(\regf[15][14] ), .S0(n1134), .S1(n1439), .Q(
        n1589) );
  MUX41X1 U2240 ( .IN1(\regf[8][14] ), .IN3(\regf[10][14] ), .IN2(
        \regf[9][14] ), .IN4(\regf[11][14] ), .S0(n1301), .S1(n1423), .Q(n1590) );
  MUX41X1 U2241 ( .IN1(\regf[4][14] ), .IN3(\regf[6][14] ), .IN2(\regf[5][14] ), .IN4(\regf[7][14] ), .S0(n1285), .S1(n1162), .Q(n1591) );
  MUX41X1 U2242 ( .IN1(n1592), .IN3(n1590), .IN2(n1591), .IN4(n1589), .S0(
        n1905), .S1(n1899), .Q(n1593) );
  MUX41X1 U2243 ( .IN1(\regf[28][15] ), .IN3(\regf[30][15] ), .IN2(
        \regf[29][15] ), .IN4(\regf[31][15] ), .S0(n1348), .S1(n1437), .Q(
        n1594) );
  MUX41X1 U2244 ( .IN1(\regf[24][15] ), .IN3(\regf[26][15] ), .IN2(
        \regf[25][15] ), .IN4(\regf[27][15] ), .S0(n1134), .S1(n1179), .Q(
        n1595) );
  MUX41X1 U2245 ( .IN1(\regf[20][15] ), .IN3(\regf[22][15] ), .IN2(
        \regf[21][15] ), .IN4(\regf[23][15] ), .S0(n1341), .S1(n1431), .Q(
        n1596) );
  MUX41X1 U2246 ( .IN1(\regf[16][15] ), .IN3(\regf[18][15] ), .IN2(
        \regf[17][15] ), .IN4(\regf[19][15] ), .S0(n1310), .S1(n1439), .Q(
        n1597) );
  MUX41X1 U2247 ( .IN1(\regf[12][15] ), .IN3(\regf[14][15] ), .IN2(
        \regf[13][15] ), .IN4(\regf[15][15] ), .S0(n1333), .S1(n1192), .Q(
        n1599) );
  MUX41X1 U2248 ( .IN1(\regf[8][15] ), .IN3(\regf[10][15] ), .IN2(
        \regf[9][15] ), .IN4(\regf[11][15] ), .S0(n1302), .S1(n1131), .Q(n1600) );
  MUX41X1 U2249 ( .IN1(\regf[4][15] ), .IN3(\regf[6][15] ), .IN2(\regf[5][15] ), .IN4(\regf[7][15] ), .S0(n1301), .S1(n1091), .Q(n1601) );
  MUX41X1 U2250 ( .IN1(n1602), .IN3(n1600), .IN2(n1601), .IN4(n1599), .S0(
        n1905), .S1(n1899), .Q(n1603) );
  MUX41X1 U2251 ( .IN1(\regf[28][16] ), .IN3(\regf[30][16] ), .IN2(
        \regf[29][16] ), .IN4(\regf[31][16] ), .S0(n1313), .S1(n1084), .Q(
        n1604) );
  MUX41X1 U2252 ( .IN1(\regf[24][16] ), .IN3(\regf[26][16] ), .IN2(
        \regf[25][16] ), .IN4(\regf[27][16] ), .S0(n1334), .S1(n1158), .Q(
        n1605) );
  MUX41X1 U2253 ( .IN1(\regf[20][16] ), .IN3(\regf[22][16] ), .IN2(
        \regf[21][16] ), .IN4(\regf[23][16] ), .S0(n1340), .S1(n1193), .Q(
        n1606) );
  MUX41X1 U2254 ( .IN1(\regf[16][16] ), .IN3(\regf[18][16] ), .IN2(
        \regf[17][16] ), .IN4(\regf[19][16] ), .S0(n1346), .S1(n1440), .Q(
        n1607) );
  MUX41X1 U2255 ( .IN1(n1607), .IN3(n1605), .IN2(n1606), .IN4(n1604), .S0(
        n1905), .S1(n1899), .Q(n1608) );
  MUX41X1 U2256 ( .IN1(\regf[12][16] ), .IN3(\regf[14][16] ), .IN2(
        \regf[13][16] ), .IN4(\regf[15][16] ), .S0(n1134), .S1(n1072), .Q(
        n1609) );
  MUX41X1 U2257 ( .IN1(\regf[8][16] ), .IN3(\regf[10][16] ), .IN2(
        \regf[9][16] ), .IN4(\regf[11][16] ), .S0(n1299), .S1(n1433), .Q(n1610) );
  MUX41X1 U2258 ( .IN1(\regf[4][16] ), .IN3(\regf[6][16] ), .IN2(\regf[5][16] ), .IN4(\regf[7][16] ), .S0(n1303), .S1(n1440), .Q(n1611) );
  MUX41X1 U2259 ( .IN1(n1612), .IN3(n1610), .IN2(n1611), .IN4(n1609), .S0(
        n1905), .S1(n1899), .Q(n1613) );
  MUX41X1 U2260 ( .IN1(\regf[28][17] ), .IN3(\regf[30][17] ), .IN2(
        \regf[29][17] ), .IN4(\regf[31][17] ), .S0(n1311), .S1(n1441), .Q(
        n1614) );
  MUX41X1 U2261 ( .IN1(\regf[24][17] ), .IN3(\regf[26][17] ), .IN2(
        \regf[25][17] ), .IN4(\regf[27][17] ), .S0(n1333), .S1(n1193), .Q(
        n1615) );
  MUX41X1 U2262 ( .IN1(\regf[16][17] ), .IN3(\regf[18][17] ), .IN2(
        \regf[17][17] ), .IN4(\regf[19][17] ), .S0(n1312), .S1(n1086), .Q(
        n1617) );
  MUX41X1 U2263 ( .IN1(\regf[12][17] ), .IN3(\regf[14][17] ), .IN2(
        \regf[13][17] ), .IN4(\regf[15][17] ), .S0(n1346), .S1(n1160), .Q(
        n1619) );
  MUX41X1 U2264 ( .IN1(\regf[8][17] ), .IN3(\regf[10][17] ), .IN2(
        \regf[9][17] ), .IN4(\regf[11][17] ), .S0(n1316), .S1(n1421), .Q(n1620) );
  MUX41X1 U2265 ( .IN1(\regf[4][17] ), .IN3(\regf[6][17] ), .IN2(\regf[5][17] ), .IN4(\regf[7][17] ), .S0(n1302), .S1(n1087), .Q(n1621) );
  MUX41X1 U2266 ( .IN1(n1622), .IN3(n1620), .IN2(n1621), .IN4(n1619), .S0(
        n1905), .S1(n1899), .Q(n1623) );
  MUX41X1 U2267 ( .IN1(\regf[28][18] ), .IN3(\regf[30][18] ), .IN2(
        \regf[29][18] ), .IN4(\regf[31][18] ), .S0(n1134), .S1(n1072), .Q(
        n1624) );
  MUX41X1 U2268 ( .IN1(\regf[24][18] ), .IN3(\regf[26][18] ), .IN2(
        \regf[25][18] ), .IN4(\regf[27][18] ), .S0(n1332), .S1(n1419), .Q(
        n1625) );
  MUX41X1 U2269 ( .IN1(\regf[16][18] ), .IN3(\regf[18][18] ), .IN2(
        \regf[17][18] ), .IN4(\regf[19][18] ), .S0(n1331), .S1(n1146), .Q(
        n1627) );
  MUX41X1 U2270 ( .IN1(n1627), .IN3(n1625), .IN2(n1626), .IN4(n1624), .S0(
        n1905), .S1(n1899), .Q(n1628) );
  MUX41X1 U2271 ( .IN1(\regf[12][18] ), .IN3(\regf[14][18] ), .IN2(
        \regf[13][18] ), .IN4(\regf[15][18] ), .S0(n1340), .S1(n1402), .Q(
        n1629) );
  MUX41X1 U2272 ( .IN1(\regf[8][18] ), .IN3(\regf[10][18] ), .IN2(
        \regf[9][18] ), .IN4(\regf[11][18] ), .S0(n1309), .S1(n1430), .Q(n1630) );
  MUX41X1 U2273 ( .IN1(\regf[4][18] ), .IN3(\regf[6][18] ), .IN2(\regf[5][18] ), .IN4(\regf[7][18] ), .S0(n1306), .S1(n1409), .Q(n1631) );
  MUX41X1 U2274 ( .IN1(n1632), .IN3(n1630), .IN2(n1631), .IN4(n1629), .S0(
        n1905), .S1(n1899), .Q(n1633) );
  MUX41X1 U2275 ( .IN1(\regf[28][19] ), .IN3(\regf[30][19] ), .IN2(
        \regf[29][19] ), .IN4(\regf[31][19] ), .S0(n1332), .S1(n1409), .Q(
        n1634) );
  MUX41X1 U2276 ( .IN1(\regf[24][19] ), .IN3(\regf[26][19] ), .IN2(
        \regf[25][19] ), .IN4(\regf[27][19] ), .S0(n1340), .S1(n1421), .Q(
        n1635) );
  MUX41X1 U2277 ( .IN1(\regf[16][19] ), .IN3(\regf[18][19] ), .IN2(
        \regf[17][19] ), .IN4(\regf[19][19] ), .S0(n1285), .S1(n1194), .Q(
        n1637) );
  MUX41X1 U2278 ( .IN1(n1637), .IN3(n1635), .IN2(n1636), .IN4(n1634), .S0(
        n1905), .S1(n1899), .Q(n1638) );
  MUX41X1 U2279 ( .IN1(\regf[8][19] ), .IN3(\regf[10][19] ), .IN2(
        \regf[9][19] ), .IN4(\regf[11][19] ), .S0(n1348), .S1(n1423), .Q(n1640) );
  MUX41X1 U2280 ( .IN1(\regf[4][19] ), .IN3(\regf[6][19] ), .IN2(\regf[5][19] ), .IN4(\regf[7][19] ), .S0(n1346), .S1(n1441), .Q(n1641) );
  MUX41X1 U2281 ( .IN1(n1642), .IN3(n1640), .IN2(n1641), .IN4(n1639), .S0(
        n1905), .S1(n1899), .Q(n1643) );
  MUX41X1 U2282 ( .IN1(\regf[28][20] ), .IN3(\regf[30][20] ), .IN2(
        \regf[29][20] ), .IN4(\regf[31][20] ), .S0(n1286), .S1(n1161), .Q(
        n1644) );
  MUX41X1 U2283 ( .IN1(\regf[24][20] ), .IN3(\regf[26][20] ), .IN2(
        \regf[25][20] ), .IN4(\regf[27][20] ), .S0(n1289), .S1(n1441), .Q(
        n1645) );
  MUX41X1 U2284 ( .IN1(\regf[20][20] ), .IN3(\regf[22][20] ), .IN2(
        \regf[21][20] ), .IN4(\regf[23][20] ), .S0(n1326), .S1(n1161), .Q(
        n1646) );
  MUX41X1 U2285 ( .IN1(\regf[16][20] ), .IN3(\regf[18][20] ), .IN2(
        \regf[17][20] ), .IN4(\regf[19][20] ), .S0(n1283), .S1(n1086), .Q(
        n1647) );
  MUX41X1 U2286 ( .IN1(n1647), .IN3(n1645), .IN2(n1646), .IN4(n1644), .S0(
        n1906), .S1(n1900), .Q(n1648) );
  MUX41X1 U2287 ( .IN1(\regf[12][20] ), .IN3(\regf[14][20] ), .IN2(
        \regf[13][20] ), .IN4(\regf[15][20] ), .S0(n1285), .S1(n1131), .Q(
        n1649) );
  MUX41X1 U2288 ( .IN1(\regf[8][20] ), .IN3(\regf[10][20] ), .IN2(
        \regf[9][20] ), .IN4(\regf[11][20] ), .S0(n1334), .S1(n1073), .Q(n1650) );
  MUX41X1 U2289 ( .IN1(\regf[4][20] ), .IN3(\regf[6][20] ), .IN2(\regf[5][20] ), .IN4(\regf[7][20] ), .S0(n1289), .S1(n1439), .Q(n1651) );
  MUX41X1 U2290 ( .IN1(n1652), .IN3(n1650), .IN2(n1651), .IN4(n1649), .S0(
        n1906), .S1(n1900), .Q(n1653) );
  MUX21X1 U2291 ( .IN1(n1653), .IN2(n1648), .S(n1910), .Q(rd_dataA[20]) );
  MUX41X1 U2292 ( .IN1(\regf[28][21] ), .IN3(\regf[30][21] ), .IN2(
        \regf[29][21] ), .IN4(\regf[31][21] ), .S0(n1333), .S1(n1428), .Q(
        n1654) );
  MUX41X1 U2293 ( .IN1(\regf[24][21] ), .IN3(\regf[26][21] ), .IN2(
        \regf[25][21] ), .IN4(\regf[27][21] ), .S0(n1290), .S1(n1131), .Q(
        n1655) );
  MUX41X1 U2294 ( .IN1(\regf[20][21] ), .IN3(\regf[22][21] ), .IN2(
        \regf[21][21] ), .IN4(\regf[23][21] ), .S0(n1287), .S1(n1436), .Q(
        n1656) );
  MUX41X1 U2295 ( .IN1(\regf[16][21] ), .IN3(\regf[18][21] ), .IN2(
        \regf[17][21] ), .IN4(\regf[19][21] ), .S0(n1346), .S1(n1180), .Q(
        n1657) );
  MUX41X1 U2296 ( .IN1(\regf[12][21] ), .IN3(\regf[14][21] ), .IN2(
        \regf[13][21] ), .IN4(\regf[15][21] ), .S0(n1290), .S1(n1151), .Q(
        n1659) );
  MUX41X1 U2297 ( .IN1(\regf[8][21] ), .IN3(\regf[10][21] ), .IN2(
        \regf[9][21] ), .IN4(\regf[11][21] ), .S0(n1295), .S1(n1192), .Q(n1660) );
  MUX41X1 U2298 ( .IN1(n1662), .IN3(n1660), .IN2(n1661), .IN4(n1659), .S0(
        n1906), .S1(n1900), .Q(n1663) );
  MUX41X1 U2299 ( .IN1(\regf[28][22] ), .IN3(\regf[30][22] ), .IN2(
        \regf[29][22] ), .IN4(\regf[31][22] ), .S0(n1288), .S1(n1127), .Q(
        n1664) );
  MUX41X1 U2300 ( .IN1(\regf[24][22] ), .IN3(\regf[26][22] ), .IN2(
        \regf[25][22] ), .IN4(\regf[27][22] ), .S0(n1291), .S1(n1437), .Q(
        n1665) );
  MUX41X1 U2301 ( .IN1(\regf[20][22] ), .IN3(\regf[22][22] ), .IN2(
        \regf[21][22] ), .IN4(\regf[23][22] ), .S0(n1290), .S1(n1177), .Q(
        n1666) );
  MUX41X1 U2302 ( .IN1(n1667), .IN3(n1665), .IN2(n1666), .IN4(n1664), .S0(
        n1906), .S1(n1900), .Q(n1668) );
  MUX41X1 U2303 ( .IN1(\regf[12][22] ), .IN3(\regf[14][22] ), .IN2(
        \regf[13][22] ), .IN4(\regf[15][22] ), .S0(n1353), .S1(n1405), .Q(
        n1669) );
  MUX41X1 U2304 ( .IN1(\regf[8][22] ), .IN3(\regf[10][22] ), .IN2(
        \regf[9][22] ), .IN4(\regf[11][22] ), .S0(n1310), .S1(n1418), .Q(n1670) );
  MUX41X1 U2305 ( .IN1(n1672), .IN3(n1670), .IN2(n1671), .IN4(n1669), .S0(
        n1906), .S1(n1900), .Q(n1673) );
  MUX41X1 U2306 ( .IN1(\regf[28][23] ), .IN3(\regf[30][23] ), .IN2(
        \regf[29][23] ), .IN4(\regf[31][23] ), .S0(n1344), .S1(n1184), .Q(
        n1674) );
  MUX41X1 U2307 ( .IN1(\regf[20][23] ), .IN3(\regf[22][23] ), .IN2(
        \regf[21][23] ), .IN4(\regf[23][23] ), .S0(n1327), .S1(n1404), .Q(
        n1676) );
  MUX41X1 U2308 ( .IN1(n1677), .IN3(n1675), .IN2(n1676), .IN4(n1674), .S0(
        n1906), .S1(n1900), .Q(n1678) );
  MUX41X1 U2309 ( .IN1(\regf[12][23] ), .IN3(\regf[14][23] ), .IN2(
        \regf[13][23] ), .IN4(\regf[15][23] ), .S0(n1283), .S1(n1150), .Q(
        n1679) );
  MUX41X1 U2310 ( .IN1(\regf[8][23] ), .IN3(\regf[10][23] ), .IN2(
        \regf[9][23] ), .IN4(\regf[11][23] ), .S0(n1296), .S1(n1398), .Q(n1680) );
  MUX41X1 U2311 ( .IN1(\regf[4][23] ), .IN3(\regf[6][23] ), .IN2(\regf[5][23] ), .IN4(\regf[7][23] ), .S0(n1348), .S1(n1079), .Q(n1681) );
  MUX41X1 U2312 ( .IN1(n1682), .IN3(n1680), .IN2(n1681), .IN4(n1679), .S0(
        n1906), .S1(n1900), .Q(n1683) );
  MUX21X1 U2313 ( .IN1(n1683), .IN2(n1678), .S(n1910), .Q(rd_dataA[23]) );
  MUX41X1 U2314 ( .IN1(\regf[28][24] ), .IN3(\regf[30][24] ), .IN2(
        \regf[29][24] ), .IN4(\regf[31][24] ), .S0(n1345), .S1(n1174), .Q(
        n1684) );
  MUX41X1 U2315 ( .IN1(\regf[24][24] ), .IN3(\regf[26][24] ), .IN2(
        \regf[25][24] ), .IN4(\regf[27][24] ), .S0(n1293), .S1(n1438), .Q(
        n1685) );
  MUX41X1 U2316 ( .IN1(\regf[20][24] ), .IN3(\regf[22][24] ), .IN2(
        \regf[21][24] ), .IN4(\regf[23][24] ), .S0(n1328), .S1(n1174), .Q(
        n1686) );
  MUX41X1 U2317 ( .IN1(\regf[16][24] ), .IN3(\regf[18][24] ), .IN2(
        \regf[17][24] ), .IN4(\regf[19][24] ), .S0(n1349), .S1(n1123), .Q(
        n1687) );
  MUX41X1 U2318 ( .IN1(n1687), .IN3(n1685), .IN2(n1686), .IN4(n1684), .S0(
        n1906), .S1(n1900), .Q(n1688) );
  MUX41X1 U2319 ( .IN1(\regf[12][24] ), .IN3(\regf[14][24] ), .IN2(
        \regf[13][24] ), .IN4(\regf[15][24] ), .S0(n1284), .S1(n1120), .Q(
        n1689) );
  MUX41X1 U2320 ( .IN1(\regf[8][24] ), .IN3(\regf[10][24] ), .IN2(
        \regf[9][24] ), .IN4(\regf[11][24] ), .S0(n1311), .S1(n1111), .Q(n1690) );
  MUX41X1 U2321 ( .IN1(\regf[4][24] ), .IN3(\regf[6][24] ), .IN2(\regf[5][24] ), .IN4(\regf[7][24] ), .S0(n1349), .S1(n1197), .Q(n1691) );
  MUX41X1 U2322 ( .IN1(n1692), .IN3(n1690), .IN2(n1691), .IN4(n1689), .S0(
        n1906), .S1(n1900), .Q(n1693) );
  MUX41X1 U2323 ( .IN1(\regf[28][25] ), .IN3(\regf[30][25] ), .IN2(
        \regf[29][25] ), .IN4(\regf[31][25] ), .S0(n1286), .S1(n1160), .Q(
        n1694) );
  MUX41X1 U2324 ( .IN1(\regf[24][25] ), .IN3(\regf[26][25] ), .IN2(
        \regf[25][25] ), .IN4(\regf[27][25] ), .S0(n1294), .S1(n1124), .Q(
        n1695) );
  MUX41X1 U2325 ( .IN1(\regf[20][25] ), .IN3(\regf[22][25] ), .IN2(
        \regf[21][25] ), .IN4(\regf[23][25] ), .S0(n1286), .S1(n1179), .Q(
        n1696) );
  MUX41X1 U2326 ( .IN1(\regf[16][25] ), .IN3(\regf[18][25] ), .IN2(
        \regf[17][25] ), .IN4(\regf[19][25] ), .S0(n1350), .S1(n1173), .Q(
        n1697) );
  MUX41X1 U2327 ( .IN1(n1697), .IN3(n1695), .IN2(n1696), .IN4(n1694), .S0(
        n1906), .S1(n1900), .Q(n1698) );
  MUX41X1 U2328 ( .IN1(\regf[12][25] ), .IN3(\regf[14][25] ), .IN2(
        \regf[13][25] ), .IN4(\regf[15][25] ), .S0(n1286), .S1(n1184), .Q(
        n1699) );
  MUX41X1 U2329 ( .IN1(\regf[8][25] ), .IN3(\regf[10][25] ), .IN2(
        \regf[9][25] ), .IN4(\regf[11][25] ), .S0(n1312), .S1(n1115), .Q(n1700) );
  MUX41X1 U2330 ( .IN1(\regf[4][25] ), .IN3(\regf[6][25] ), .IN2(\regf[5][25] ), .IN4(\regf[7][25] ), .S0(n1350), .S1(n1193), .Q(n1701) );
  MUX41X1 U2331 ( .IN1(n1702), .IN3(n1700), .IN2(n1701), .IN4(n1699), .S0(
        n1906), .S1(n1900), .Q(n1703) );
  MUX41X1 U2332 ( .IN1(\regf[28][26] ), .IN3(\regf[30][26] ), .IN2(
        \regf[29][26] ), .IN4(\regf[31][26] ), .S0(n1346), .S1(n1129), .Q(
        n1704) );
  MUX41X1 U2333 ( .IN1(\regf[24][26] ), .IN3(\regf[26][26] ), .IN2(
        \regf[25][26] ), .IN4(\regf[27][26] ), .S0(n1295), .S1(n1075), .Q(
        n1705) );
  MUX41X1 U2334 ( .IN1(\regf[20][26] ), .IN3(\regf[22][26] ), .IN2(
        \regf[21][26] ), .IN4(\regf[23][26] ), .S0(n1353), .S1(n1185), .Q(
        n1706) );
  MUX41X1 U2335 ( .IN1(n1707), .IN3(n1705), .IN2(n1706), .IN4(n1704), .S0(
        n1907), .S1(n1901), .Q(n1708) );
  MUX41X1 U2336 ( .IN1(\regf[12][26] ), .IN3(\regf[14][26] ), .IN2(
        \regf[13][26] ), .IN4(\regf[15][26] ), .S0(n1287), .S1(n1443), .Q(
        n1709) );
  MUX41X1 U2337 ( .IN1(\regf[8][26] ), .IN3(\regf[10][26] ), .IN2(
        \regf[9][26] ), .IN4(\regf[11][26] ), .S0(n1313), .S1(n1128), .Q(n1710) );
  MUX41X1 U2338 ( .IN1(n1712), .IN3(n1710), .IN2(n1711), .IN4(n1709), .S0(
        n1907), .S1(n1901), .Q(n1713) );
  MUX41X1 U2339 ( .IN1(\regf[28][27] ), .IN3(\regf[30][27] ), .IN2(
        \regf[29][27] ), .IN4(\regf[31][27] ), .S0(n1289), .S1(n1437), .Q(
        n1714) );
  MUX41X1 U2340 ( .IN1(\regf[24][27] ), .IN3(\regf[26][27] ), .IN2(
        \regf[25][27] ), .IN4(\regf[27][27] ), .S0(n1296), .S1(n1081), .Q(
        n1715) );
  MUX41X1 U2341 ( .IN1(\regf[20][27] ), .IN3(\regf[22][27] ), .IN2(
        \regf[21][27] ), .IN4(\regf[23][27] ), .S0(n1329), .S1(n1124), .Q(
        n1716) );
  MUX41X1 U2342 ( .IN1(n1717), .IN3(n1715), .IN2(n1716), .IN4(n1714), .S0(
        n1907), .S1(n1901), .Q(n1718) );
  MUX41X1 U2343 ( .IN1(\regf[12][27] ), .IN3(\regf[14][27] ), .IN2(
        \regf[13][27] ), .IN4(\regf[15][27] ), .S0(n1288), .S1(n1091), .Q(
        n1719) );
  MUX41X1 U2344 ( .IN1(\regf[8][27] ), .IN3(\regf[10][27] ), .IN2(
        \regf[9][27] ), .IN4(\regf[11][27] ), .S0(n1134), .S1(n1172), .Q(n1720) );
  MUX21X1 U2345 ( .IN1(n1723), .IN2(n1718), .S(n1910), .Q(rd_dataA[27]) );
  MUX41X1 U2346 ( .IN1(\regf[28][28] ), .IN3(\regf[30][28] ), .IN2(
        \regf[29][28] ), .IN4(\regf[31][28] ), .S0(n1284), .S1(n1121), .Q(
        n1724) );
  MUX41X1 U2347 ( .IN1(\regf[24][28] ), .IN3(\regf[26][28] ), .IN2(
        \regf[25][28] ), .IN4(\regf[27][28] ), .S0(n1297), .S1(n1436), .Q(
        n1725) );
  MUX41X1 U2348 ( .IN1(\regf[20][28] ), .IN3(\regf[22][28] ), .IN2(
        \regf[21][28] ), .IN4(\regf[23][28] ), .S0(n1283), .S1(n1080), .Q(
        n1726) );
  MUX41X1 U2349 ( .IN1(\regf[16][28] ), .IN3(\regf[18][28] ), .IN2(
        \regf[17][28] ), .IN4(\regf[19][28] ), .S0(n1285), .S1(n1429), .Q(
        n1727) );
  MUX41X1 U2350 ( .IN1(n1727), .IN3(n1725), .IN2(n1726), .IN4(n1724), .S0(
        n1907), .S1(n1901), .Q(n1728) );
  MUX41X1 U2351 ( .IN1(\regf[12][28] ), .IN3(\regf[14][28] ), .IN2(
        \regf[13][28] ), .IN4(\regf[15][28] ), .S0(n1289), .S1(n1115), .Q(
        n1729) );
  MUX41X1 U2352 ( .IN1(\regf[8][28] ), .IN3(\regf[10][28] ), .IN2(
        \regf[9][28] ), .IN4(\regf[11][28] ), .S0(n1314), .S1(n1410), .Q(n1730) );
  MUX41X1 U2353 ( .IN1(\regf[4][28] ), .IN3(\regf[6][28] ), .IN2(\regf[5][28] ), .IN4(\regf[7][28] ), .S0(n1288), .S1(n1149), .Q(n1731) );
  MUX41X1 U2354 ( .IN1(n1732), .IN3(n1730), .IN2(n1731), .IN4(n1729), .S0(
        n1907), .S1(n1901), .Q(n1733) );
  MUX41X1 U2355 ( .IN1(\regf[24][29] ), .IN3(\regf[26][29] ), .IN2(
        \regf[25][29] ), .IN4(\regf[27][29] ), .S0(n1298), .S1(n1196), .Q(
        n1735) );
  MUX41X1 U2356 ( .IN1(\regf[20][29] ), .IN3(\regf[22][29] ), .IN2(
        \regf[21][29] ), .IN4(\regf[23][29] ), .S0(n1330), .S1(n1178), .Q(
        n1736) );
  MUX41X1 U2357 ( .IN1(\regf[16][29] ), .IN3(\regf[18][29] ), .IN2(
        \regf[17][29] ), .IN4(\regf[19][29] ), .S0(n1353), .S1(n1162), .Q(
        n1737) );
  MUX41X1 U2358 ( .IN1(\regf[12][29] ), .IN3(\regf[14][29] ), .IN2(
        \regf[13][29] ), .IN4(\regf[15][29] ), .S0(n1290), .S1(n1441), .Q(
        n1739) );
  MUX41X1 U2359 ( .IN1(\regf[8][29] ), .IN3(\regf[10][29] ), .IN2(
        \regf[9][29] ), .IN4(\regf[11][29] ), .S0(n1315), .S1(n1419), .Q(n1740) );
  MUX41X1 U2360 ( .IN1(\regf[4][29] ), .IN3(\regf[6][29] ), .IN2(\regf[5][29] ), .IN4(\regf[7][29] ), .S0(n1315), .S1(n1114), .Q(n1741) );
  MUX41X1 U2361 ( .IN1(n1742), .IN3(n1740), .IN2(n1741), .IN4(n1739), .S0(
        n1907), .S1(n1901), .Q(n1743) );
  MUX41X1 U2362 ( .IN1(\regf[28][30] ), .IN3(\regf[30][30] ), .IN2(
        \regf[29][30] ), .IN4(\regf[31][30] ), .S0(n1290), .S1(n1074), .Q(
        n1744) );
  MUX41X1 U2363 ( .IN1(\regf[24][30] ), .IN3(\regf[26][30] ), .IN2(
        \regf[25][30] ), .IN4(\regf[27][30] ), .S0(n1283), .S1(n1076), .Q(
        n1745) );
  MUX41X1 U2364 ( .IN1(n1747), .IN3(n1745), .IN2(n1746), .IN4(n1744), .S0(
        n1907), .S1(n1901), .Q(n1748) );
  MUX41X1 U2365 ( .IN1(\regf[8][30] ), .IN3(\regf[10][30] ), .IN2(
        \regf[9][30] ), .IN4(\regf[11][30] ), .S0(n1291), .S1(n1440), .Q(n1750) );
  MUX41X1 U2366 ( .IN1(\regf[4][30] ), .IN3(\regf[6][30] ), .IN2(\regf[5][30] ), .IN4(\regf[7][30] ), .S0(n1342), .S1(n1127), .Q(n1751) );
  MUX41X1 U2367 ( .IN1(n1752), .IN3(n1750), .IN2(n1751), .IN4(n1749), .S0(
        n1907), .S1(n1901), .Q(n1753) );
  MUX41X1 U2368 ( .IN1(\regf[28][31] ), .IN3(\regf[30][31] ), .IN2(
        \regf[29][31] ), .IN4(\regf[31][31] ), .S0(n1283), .S1(n1418), .Q(
        n1754) );
  MUX41X1 U2369 ( .IN1(\regf[24][31] ), .IN3(\regf[26][31] ), .IN2(
        \regf[25][31] ), .IN4(\regf[27][31] ), .S0(n1284), .S1(n1197), .Q(
        n1755) );
  MUX41X1 U2370 ( .IN1(\regf[20][31] ), .IN3(\regf[22][31] ), .IN2(
        \regf[21][31] ), .IN4(\regf[23][31] ), .S0(n1325), .S1(n1079), .Q(
        n1756) );
  MUX41X1 U2371 ( .IN1(n1757), .IN3(n1755), .IN2(n1756), .IN4(n1754), .S0(
        n1907), .S1(n1901), .Q(n1758) );
  MUX41X1 U2372 ( .IN1(\regf[8][31] ), .IN3(\regf[10][31] ), .IN2(
        \regf[9][31] ), .IN4(\regf[11][31] ), .S0(n1292), .S1(n1076), .Q(n1760) );
  MUX41X1 U2373 ( .IN1(n1762), .IN3(n1760), .IN2(n1761), .IN4(n1759), .S0(
        n1907), .S1(n1901), .Q(n1763) );
  MUX21X1 U2374 ( .IN1(n1764), .IN2(n1765), .S(n1291), .Q(n1767) );
  MUX21X1 U2375 ( .IN1(n1768), .IN2(n1769), .S(n1313), .Q(n1771) );
  MUX21X1 U2376 ( .IN1(n1772), .IN2(n1773), .S(n1292), .Q(n1775) );
  MUX21X1 U2377 ( .IN1(n1776), .IN2(n1777), .S(n1293), .Q(n1779) );
  MUX21X1 U2378 ( .IN1(n1784), .IN2(n1785), .S(n1294), .Q(n1787) );
  MUX21X1 U2379 ( .IN1(n1788), .IN2(n1789), .S(n1295), .Q(n1791) );
  MUX21X1 U2380 ( .IN1(n1792), .IN2(n1793), .S(n1316), .Q(n1795) );
  MUX21X1 U2381 ( .IN1(n1800), .IN2(n1801), .S(n1297), .Q(n1803) );
  MUX21X1 U2382 ( .IN1(n1804), .IN2(n1805), .S(n1318), .Q(n1807) );
  MUX21X1 U2383 ( .IN1(n1808), .IN2(n1809), .S(n1298), .Q(n1811) );
  MUX21X1 U2384 ( .IN1(n1820), .IN2(n1821), .S(n1310), .Q(n1823) );
  MUX21X1 U2385 ( .IN1(n1824), .IN2(n1825), .S(n1311), .Q(n1827) );
  MUX21X1 U2386 ( .IN1(n1828), .IN2(n1829), .S(n1300), .Q(n1831) );
  MUX21X1 U2387 ( .IN1(n1832), .IN2(n1833), .S(n1312), .Q(n1835) );
  MUX21X1 U2388 ( .IN1(n1836), .IN2(n1837), .S(n1310), .Q(n1839) );
  NAND3X0 U2389 ( .IN1(\regf[3][13] ), .IN2(n1289), .IN3(n1195), .QN(n1838) );
  MUX21X1 U2390 ( .IN1(n1840), .IN2(n1841), .S(n1302), .Q(n1843) );
  MUX21X1 U2391 ( .IN1(n1844), .IN2(n1845), .S(n1315), .Q(n1847) );
  MUX21X1 U2392 ( .IN1(n1848), .IN2(n1849), .S(n1317), .Q(n1851) );
  NAND3X0 U2393 ( .IN1(\regf[3][10] ), .IN2(n1295), .IN3(n1172), .QN(n1850) );
  MUX21X1 U2394 ( .IN1(n1852), .IN2(n1853), .S(n1304), .Q(n1855) );
  MUX21X1 U2395 ( .IN1(n1856), .IN2(n1857), .S(n1299), .Q(n1859) );
  MUX21X1 U2396 ( .IN1(n1860), .IN2(n1861), .S(n1301), .Q(n1863) );
  MUX21X1 U2397 ( .IN1(n1864), .IN2(n1865), .S(n1306), .Q(n1867) );
  MUX21X1 U2398 ( .IN1(n1876), .IN2(n1877), .S(n1308), .Q(n1879) );
  MUX21X1 U2399 ( .IN1(n1880), .IN2(n1881), .S(n1307), .Q(n1883) );
  NAND3X0 U2400 ( .IN1(\regf[3][1] ), .IN2(n1294), .IN3(n1162), .QN(n1886) );
  MUX21X1 U2401 ( .IN1(n1888), .IN2(n1889), .S(n1308), .Q(n1891) );
  NAND3X0 U2402 ( .IN1(\regf[3][0] ), .IN2(n1289), .IN3(n1434), .QN(n1890) );
  INVX0 U2403 ( .INP(N11), .ZN(n1892) );
  DELLN1X2 U2404 ( .INP(n1892), .Z(n1893) );
  DELLN1X2 U2405 ( .INP(N12), .Z(n1895) );
  DELLN1X2 U2406 ( .INP(N13), .Z(n1897) );
  DELLN1X2 U2407 ( .INP(N13), .Z(n1898) );
  DELLN1X2 U2408 ( .INP(N13), .Z(n1899) );
  DELLN1X2 U2409 ( .INP(N13), .Z(n1900) );
  DELLN1X2 U2410 ( .INP(N13), .Z(n1901) );
  DELLN1X2 U2411 ( .INP(N15), .Z(n1910) );
  DELLN1X2 U2412 ( .INP(N14), .Z(n1906) );
  DELLN1X2 U2413 ( .INP(N14), .Z(n1907) );
  MUX41X1 U2414 ( .IN1(\regf[28][0] ), .IN3(\regf[30][0] ), .IN2(\regf[29][0] ), .IN4(\regf[31][0] ), .S0(n1208), .S1(n1191), .Q(n1911) );
  MUX41X1 U2415 ( .IN1(\regf[24][0] ), .IN3(\regf[26][0] ), .IN2(\regf[25][0] ), .IN4(\regf[27][0] ), .S0(n1209), .S1(n1385), .Q(n1912) );
  MUX41X1 U2416 ( .IN1(\regf[20][0] ), .IN3(\regf[22][0] ), .IN2(\regf[21][0] ), .IN4(\regf[23][0] ), .S0(n1270), .S1(n1135), .Q(n1913) );
  MUX41X1 U2417 ( .IN1(\regf[16][0] ), .IN3(\regf[18][0] ), .IN2(\regf[17][0] ), .IN4(\regf[19][0] ), .S0(n1265), .S1(n1392), .Q(n1914) );
  MUX41X1 U2418 ( .IN1(n1914), .IN3(n1912), .IN2(n1913), .IN4(n1911), .S0(
        n2374), .S1(n2368), .Q(n1915) );
  MUX41X1 U2419 ( .IN1(\regf[12][0] ), .IN3(\regf[14][0] ), .IN2(\regf[13][0] ), .IN4(\regf[15][0] ), .S0(n1271), .S1(n1390), .Q(n1916) );
  MUX41X1 U2420 ( .IN1(\regf[8][0] ), .IN3(\regf[10][0] ), .IN2(\regf[9][0] ), 
        .IN4(\regf[11][0] ), .S0(n1214), .S1(n1365), .Q(n1917) );
  MUX41X1 U2421 ( .IN1(\regf[4][0] ), .IN3(\regf[6][0] ), .IN2(\regf[5][0] ), 
        .IN4(\regf[7][0] ), .S0(n1267), .S1(n1166), .Q(n1918) );
  MUX41X1 U2422 ( .IN1(n1919), .IN3(n1917), .IN2(n1918), .IN4(n1916), .S0(
        n2374), .S1(n2368), .Q(n1920) );
  MUX41X1 U2423 ( .IN1(\regf[28][1] ), .IN3(\regf[30][1] ), .IN2(\regf[29][1] ), .IN4(\regf[31][1] ), .S0(n1266), .S1(n1135), .Q(n1921) );
  MUX41X1 U2424 ( .IN1(\regf[24][1] ), .IN3(\regf[26][1] ), .IN2(\regf[25][1] ), .IN4(\regf[27][1] ), .S0(n1206), .S1(n1374), .Q(n1922) );
  MUX41X1 U2425 ( .IN1(\regf[20][1] ), .IN3(\regf[22][1] ), .IN2(\regf[21][1] ), .IN4(\regf[23][1] ), .S0(n1271), .S1(n1387), .Q(n1923) );
  MUX41X1 U2426 ( .IN1(\regf[16][1] ), .IN3(\regf[18][1] ), .IN2(\regf[17][1] ), .IN4(\regf[19][1] ), .S0(n1210), .S1(n1372), .Q(n1924) );
  MUX41X1 U2427 ( .IN1(n1924), .IN3(n1922), .IN2(n1923), .IN4(n1921), .S0(
        n2374), .S1(n2368), .Q(n1925) );
  MUX41X1 U2428 ( .IN1(\regf[12][1] ), .IN3(\regf[14][1] ), .IN2(\regf[13][1] ), .IN4(\regf[15][1] ), .S0(n1272), .S1(n1383), .Q(n1926) );
  MUX41X1 U2429 ( .IN1(\regf[8][1] ), .IN3(\regf[10][1] ), .IN2(\regf[9][1] ), 
        .IN4(\regf[11][1] ), .S0(n1215), .S1(n1366), .Q(n1927) );
  MUX41X1 U2430 ( .IN1(\regf[4][1] ), .IN3(\regf[6][1] ), .IN2(\regf[5][1] ), 
        .IN4(\regf[7][1] ), .S0(n1266), .S1(n1170), .Q(n1928) );
  MUX41X1 U2431 ( .IN1(n1929), .IN3(n1927), .IN2(n1928), .IN4(n1926), .S0(
        n2374), .S1(n2368), .Q(n1930) );
  MUX21X1 U2432 ( .IN1(n1930), .IN2(n1925), .S(n2380), .Q(rd_dataB[1]) );
  MUX41X1 U2433 ( .IN1(\regf[28][2] ), .IN3(\regf[30][2] ), .IN2(\regf[29][2] ), .IN4(\regf[31][2] ), .S0(n1205), .S1(n1354), .Q(n1931) );
  MUX41X1 U2434 ( .IN1(\regf[24][2] ), .IN3(\regf[26][2] ), .IN2(\regf[25][2] ), .IN4(\regf[27][2] ), .S0(n1207), .S1(n1147), .Q(n1932) );
  MUX41X1 U2435 ( .IN1(\regf[20][2] ), .IN3(\regf[22][2] ), .IN2(\regf[21][2] ), .IN4(\regf[23][2] ), .S0(n1272), .S1(n1377), .Q(n1933) );
  MUX41X1 U2436 ( .IN1(\regf[16][2] ), .IN3(\regf[18][2] ), .IN2(\regf[17][2] ), .IN4(\regf[19][2] ), .S0(n1267), .S1(n1168), .Q(n1934) );
  MUX41X1 U2437 ( .IN1(n1934), .IN3(n1932), .IN2(n1933), .IN4(n1931), .S0(
        n2375), .S1(n2369), .Q(n1935) );
  MUX41X1 U2438 ( .IN1(\regf[12][2] ), .IN3(\regf[14][2] ), .IN2(\regf[13][2] ), .IN4(\regf[15][2] ), .S0(n1273), .S1(n1377), .Q(n1936) );
  MUX41X1 U2439 ( .IN1(\regf[8][2] ), .IN3(\regf[10][2] ), .IN2(\regf[9][2] ), 
        .IN4(\regf[11][2] ), .S0(n1267), .S1(n1096), .Q(n1937) );
  MUX41X1 U2440 ( .IN1(\regf[4][2] ), .IN3(\regf[6][2] ), .IN2(\regf[5][2] ), 
        .IN4(\regf[7][2] ), .S0(n1220), .S1(n1394), .Q(n1938) );
  MUX41X1 U2441 ( .IN1(n1939), .IN3(n1937), .IN2(n1938), .IN4(n1936), .S0(
        n2375), .S1(n2369), .Q(n1940) );
  MUX41X1 U2442 ( .IN1(\regf[28][3] ), .IN3(\regf[30][3] ), .IN2(\regf[29][3] ), .IN4(\regf[31][3] ), .S0(n1204), .S1(n1092), .Q(n1941) );
  MUX41X1 U2443 ( .IN1(\regf[24][3] ), .IN3(\regf[26][3] ), .IN2(\regf[25][3] ), .IN4(\regf[27][3] ), .S0(n1262), .S1(n1382), .Q(n1942) );
  MUX41X1 U2444 ( .IN1(\regf[20][3] ), .IN3(\regf[22][3] ), .IN2(\regf[21][3] ), .IN4(\regf[23][3] ), .S0(n1260), .S1(n1385), .Q(n1943) );
  MUX41X1 U2445 ( .IN1(\regf[16][3] ), .IN3(\regf[18][3] ), .IN2(\regf[17][3] ), .IN4(\regf[19][3] ), .S0(n1255), .S1(n1393), .Q(n1944) );
  MUX41X1 U2446 ( .IN1(n1944), .IN3(n1942), .IN2(n1943), .IN4(n1941), .S0(
        n2375), .S1(n2369), .Q(n1945) );
  MUX41X1 U2447 ( .IN1(\regf[12][3] ), .IN3(\regf[14][3] ), .IN2(\regf[13][3] ), .IN4(\regf[15][3] ), .S0(n1264), .S1(n1376), .Q(n1946) );
  MUX41X1 U2448 ( .IN1(\regf[8][3] ), .IN3(\regf[10][3] ), .IN2(\regf[9][3] ), 
        .IN4(\regf[11][3] ), .S0(n1237), .S1(n1095), .Q(n1947) );
  MUX41X1 U2449 ( .IN1(\regf[4][3] ), .IN3(\regf[6][3] ), .IN2(\regf[5][3] ), 
        .IN4(\regf[7][3] ), .S0(n1221), .S1(n1382), .Q(n1948) );
  MUX41X1 U2450 ( .IN1(\regf[28][4] ), .IN3(\regf[30][4] ), .IN2(\regf[29][4] ), .IN4(\regf[31][4] ), .S0(n1258), .S1(n1157), .Q(n1951) );
  MUX41X1 U2451 ( .IN1(\regf[24][4] ), .IN3(\regf[26][4] ), .IN2(\regf[25][4] ), .IN4(\regf[27][4] ), .S0(n1264), .S1(n1364), .Q(n1952) );
  MUX41X1 U2452 ( .IN1(\regf[20][4] ), .IN3(\regf[22][4] ), .IN2(\regf[21][4] ), .IN4(\regf[23][4] ), .S0(n1257), .S1(n1089), .Q(n1953) );
  MUX41X1 U2453 ( .IN1(\regf[16][4] ), .IN3(\regf[18][4] ), .IN2(\regf[17][4] ), .IN4(\regf[19][4] ), .S0(n1256), .S1(n1364), .Q(n1954) );
  MUX41X1 U2454 ( .IN1(n1954), .IN3(n1952), .IN2(n1953), .IN4(n1951), .S0(
        n2375), .S1(n2369), .Q(n1955) );
  MUX41X1 U2455 ( .IN1(\regf[12][4] ), .IN3(\regf[14][4] ), .IN2(\regf[13][4] ), .IN4(\regf[15][4] ), .S0(n1261), .S1(n1169), .Q(n1956) );
  MUX41X1 U2456 ( .IN1(\regf[8][4] ), .IN3(\regf[10][4] ), .IN2(\regf[9][4] ), 
        .IN4(\regf[11][4] ), .S0(n1238), .S1(n1359), .Q(n1957) );
  MUX41X1 U2457 ( .IN1(\regf[4][4] ), .IN3(\regf[6][4] ), .IN2(\regf[5][4] ), 
        .IN4(\regf[7][4] ), .S0(n1211), .S1(n1155), .Q(n1958) );
  MUX41X1 U2458 ( .IN1(n1959), .IN3(n1957), .IN2(n1958), .IN4(n1956), .S0(
        n2375), .S1(n2369), .Q(n1960) );
  MUX41X1 U2459 ( .IN1(\regf[28][5] ), .IN3(\regf[30][5] ), .IN2(\regf[29][5] ), .IN4(\regf[31][5] ), .S0(n1246), .S1(n1094), .Q(n1961) );
  MUX41X1 U2460 ( .IN1(\regf[24][5] ), .IN3(\regf[26][5] ), .IN2(\regf[25][5] ), .IN4(\regf[27][5] ), .S0(n1209), .S1(n1365), .Q(n1962) );
  MUX41X1 U2461 ( .IN1(\regf[20][5] ), .IN3(\regf[22][5] ), .IN2(\regf[21][5] ), .IN4(\regf[23][5] ), .S0(n1209), .S1(n1113), .Q(n1963) );
  MUX41X1 U2462 ( .IN1(\regf[16][5] ), .IN3(\regf[18][5] ), .IN2(\regf[17][5] ), .IN4(\regf[19][5] ), .S0(n1250), .S1(n1355), .Q(n1964) );
  MUX41X1 U2463 ( .IN1(n1964), .IN3(n1962), .IN2(n1963), .IN4(n1961), .S0(
        n2375), .S1(n2369), .Q(n1965) );
  MUX41X1 U2464 ( .IN1(\regf[12][5] ), .IN3(\regf[14][5] ), .IN2(\regf[13][5] ), .IN4(\regf[15][5] ), .S0(n1204), .S1(n1145), .Q(n1966) );
  MUX41X1 U2465 ( .IN1(\regf[8][5] ), .IN3(\regf[10][5] ), .IN2(\regf[9][5] ), 
        .IN4(\regf[11][5] ), .S0(n1228), .S1(n1392), .Q(n1967) );
  MUX41X1 U2466 ( .IN1(\regf[4][5] ), .IN3(\regf[6][5] ), .IN2(\regf[5][5] ), 
        .IN4(\regf[7][5] ), .S0(n1225), .S1(n1363), .Q(n1968) );
  MUX21X1 U2467 ( .IN1(n1970), .IN2(n1965), .S(n2380), .Q(rd_dataB[5]) );
  MUX41X1 U2468 ( .IN1(\regf[28][6] ), .IN3(\regf[30][6] ), .IN2(\regf[29][6] ), .IN4(\regf[31][6] ), .S0(n1248), .S1(n1372), .Q(n1971) );
  MUX41X1 U2469 ( .IN1(\regf[24][6] ), .IN3(\regf[26][6] ), .IN2(\regf[25][6] ), .IN4(\regf[27][6] ), .S0(n1259), .S1(n1376), .Q(n1972) );
  MUX41X1 U2470 ( .IN1(\regf[20][6] ), .IN3(\regf[22][6] ), .IN2(\regf[21][6] ), .IN4(\regf[23][6] ), .S0(n1267), .S1(n1354), .Q(n1973) );
  MUX41X1 U2471 ( .IN1(\regf[16][6] ), .IN3(\regf[18][6] ), .IN2(\regf[17][6] ), .IN4(\regf[19][6] ), .S0(n1251), .S1(n1382), .Q(n1974) );
  MUX41X1 U2472 ( .IN1(n1974), .IN3(n1972), .IN2(n1973), .IN4(n1971), .S0(
        n2375), .S1(n2369), .Q(n1975) );
  MUX41X1 U2473 ( .IN1(\regf[12][6] ), .IN3(\regf[14][6] ), .IN2(\regf[13][6] ), .IN4(\regf[15][6] ), .S0(n1260), .S1(n1387), .Q(n1976) );
  MUX41X1 U2474 ( .IN1(\regf[8][6] ), .IN3(\regf[10][6] ), .IN2(\regf[9][6] ), 
        .IN4(\regf[11][6] ), .S0(n1229), .S1(n1391), .Q(n1977) );
  MUX41X1 U2475 ( .IN1(\regf[4][6] ), .IN3(\regf[6][6] ), .IN2(\regf[5][6] ), 
        .IN4(\regf[7][6] ), .S0(n1226), .S1(n1168), .Q(n1978) );
  MUX21X1 U2476 ( .IN1(n1980), .IN2(n1975), .S(n2380), .Q(rd_dataB[6]) );
  MUX41X1 U2477 ( .IN1(\regf[28][7] ), .IN3(\regf[30][7] ), .IN2(\regf[29][7] ), .IN4(\regf[31][7] ), .S0(n1238), .S1(n1394), .Q(n1981) );
  MUX41X1 U2478 ( .IN1(\regf[24][7] ), .IN3(\regf[26][7] ), .IN2(\regf[25][7] ), .IN4(\regf[27][7] ), .S0(n1216), .S1(n1164), .Q(n1982) );
  MUX41X1 U2479 ( .IN1(\regf[20][7] ), .IN3(\regf[22][7] ), .IN2(\regf[21][7] ), .IN4(\regf[23][7] ), .S0(n1266), .S1(n1137), .Q(n1983) );
  MUX41X1 U2480 ( .IN1(\regf[16][7] ), .IN3(\regf[18][7] ), .IN2(\regf[17][7] ), .IN4(\regf[19][7] ), .S0(n1204), .S1(n1374), .Q(n1984) );
  MUX41X1 U2481 ( .IN1(\regf[12][7] ), .IN3(\regf[14][7] ), .IN2(\regf[13][7] ), .IN4(\regf[15][7] ), .S0(n1259), .S1(n1071), .Q(n1986) );
  MUX41X1 U2482 ( .IN1(\regf[8][7] ), .IN3(\regf[10][7] ), .IN2(\regf[9][7] ), 
        .IN4(\regf[11][7] ), .S0(n1226), .S1(n1113), .Q(n1987) );
  MUX41X1 U2483 ( .IN1(\regf[4][7] ), .IN3(\regf[6][7] ), .IN2(\regf[5][7] ), 
        .IN4(\regf[7][7] ), .S0(n1209), .S1(n1382), .Q(n1988) );
  MUX41X1 U2484 ( .IN1(n1989), .IN3(n1987), .IN2(n1988), .IN4(n1986), .S0(
        n2375), .S1(n2369), .Q(n1990) );
  MUX41X1 U2485 ( .IN1(\regf[28][8] ), .IN3(\regf[30][8] ), .IN2(\regf[29][8] ), .IN4(\regf[31][8] ), .S0(n1126), .S1(n1154), .Q(n1991) );
  MUX41X1 U2486 ( .IN1(\regf[24][8] ), .IN3(\regf[26][8] ), .IN2(\regf[25][8] ), .IN4(\regf[27][8] ), .S0(n1208), .S1(n1377), .Q(n1992) );
  MUX41X1 U2487 ( .IN1(\regf[20][8] ), .IN3(\regf[22][8] ), .IN2(\regf[21][8] ), .IN4(\regf[23][8] ), .S0(n1266), .S1(n1383), .Q(n1993) );
  MUX41X1 U2488 ( .IN1(\regf[16][8] ), .IN3(\regf[18][8] ), .IN2(\regf[17][8] ), .IN4(\regf[19][8] ), .S0(n1207), .S1(n1363), .Q(n1994) );
  MUX41X1 U2489 ( .IN1(\regf[12][8] ), .IN3(\regf[14][8] ), .IN2(\regf[13][8] ), .IN4(\regf[15][8] ), .S0(n1257), .S1(n1376), .Q(n1996) );
  MUX41X1 U2490 ( .IN1(\regf[8][8] ), .IN3(\regf[10][8] ), .IN2(\regf[9][8] ), 
        .IN4(\regf[11][8] ), .S0(n1227), .S1(n1112), .Q(n1997) );
  MUX41X1 U2491 ( .IN1(\regf[4][8] ), .IN3(\regf[6][8] ), .IN2(\regf[5][8] ), 
        .IN4(\regf[7][8] ), .S0(n1210), .S1(n1391), .Q(n1998) );
  MUX41X1 U2492 ( .IN1(n1999), .IN3(n1997), .IN2(n1998), .IN4(n1996), .S0(
        n2376), .S1(n2370), .Q(n2000) );
  MUX41X1 U2493 ( .IN1(\regf[28][9] ), .IN3(\regf[30][9] ), .IN2(\regf[29][9] ), .IN4(\regf[31][9] ), .S0(n1245), .S1(n1355), .Q(n2001) );
  MUX41X1 U2494 ( .IN1(\regf[24][9] ), .IN3(\regf[26][9] ), .IN2(\regf[25][9] ), .IN4(\regf[27][9] ), .S0(n1248), .S1(n1181), .Q(n2002) );
  MUX41X1 U2495 ( .IN1(\regf[20][9] ), .IN3(\regf[22][9] ), .IN2(\regf[21][9] ), .IN4(\regf[23][9] ), .S0(n1206), .S1(n1387), .Q(n2003) );
  MUX41X1 U2496 ( .IN1(\regf[16][9] ), .IN3(\regf[18][9] ), .IN2(\regf[17][9] ), .IN4(\regf[19][9] ), .S0(n1228), .S1(n1145), .Q(n2004) );
  MUX41X1 U2497 ( .IN1(\regf[12][9] ), .IN3(\regf[14][9] ), .IN2(\regf[13][9] ), .IN4(\regf[15][9] ), .S0(n1248), .S1(n1396), .Q(n2006) );
  MUX41X1 U2498 ( .IN1(\regf[8][9] ), .IN3(\regf[10][9] ), .IN2(\regf[9][9] ), 
        .IN4(\regf[11][9] ), .S0(n1218), .S1(n1377), .Q(n2007) );
  MUX41X1 U2499 ( .IN1(\regf[4][9] ), .IN3(\regf[6][9] ), .IN2(\regf[5][9] ), 
        .IN4(\regf[7][9] ), .S0(n1206), .S1(n1093), .Q(n2008) );
  MUX41X1 U2500 ( .IN1(n2009), .IN3(n2007), .IN2(n2008), .IN4(n2006), .S0(
        n2376), .S1(n2370), .Q(n2010) );
  MUX41X1 U2501 ( .IN1(\regf[28][10] ), .IN3(\regf[30][10] ), .IN2(
        \regf[29][10] ), .IN4(\regf[31][10] ), .S0(n1229), .S1(n1390), .Q(
        n2011) );
  MUX41X1 U2502 ( .IN1(\regf[24][10] ), .IN3(\regf[26][10] ), .IN2(
        \regf[25][10] ), .IN4(\regf[27][10] ), .S0(n1253), .S1(n1104), .Q(
        n2012) );
  MUX41X1 U2503 ( .IN1(\regf[20][10] ), .IN3(\regf[22][10] ), .IN2(
        \regf[21][10] ), .IN4(\regf[23][10] ), .S0(n1259), .S1(n1383), .Q(
        n2013) );
  MUX41X1 U2504 ( .IN1(\regf[16][10] ), .IN3(\regf[18][10] ), .IN2(
        \regf[17][10] ), .IN4(\regf[19][10] ), .S0(n1267), .S1(n1385), .Q(
        n2014) );
  MUX41X1 U2505 ( .IN1(n2014), .IN3(n2012), .IN2(n2013), .IN4(n2011), .S0(
        n2376), .S1(n2370), .Q(n2015) );
  MUX41X1 U2506 ( .IN1(\regf[12][10] ), .IN3(\regf[14][10] ), .IN2(
        \regf[13][10] ), .IN4(\regf[15][10] ), .S0(n1250), .S1(n1110), .Q(
        n2016) );
  MUX41X1 U2507 ( .IN1(\regf[8][10] ), .IN3(\regf[10][10] ), .IN2(
        \regf[9][10] ), .IN4(\regf[11][10] ), .S0(n1219), .S1(n1394), .Q(n2017) );
  MUX41X1 U2508 ( .IN1(\regf[4][10] ), .IN3(\regf[6][10] ), .IN2(\regf[5][10] ), .IN4(\regf[7][10] ), .S0(n1204), .S1(n1088), .Q(n2018) );
  MUX41X1 U2509 ( .IN1(n2019), .IN3(n2017), .IN2(n2018), .IN4(n2016), .S0(
        n2376), .S1(n2370), .Q(n2020) );
  MUX41X1 U2510 ( .IN1(\regf[28][11] ), .IN3(\regf[30][11] ), .IN2(
        \regf[29][11] ), .IN4(\regf[31][11] ), .S0(n1230), .S1(n1355), .Q(
        n2021) );
  MUX41X1 U2511 ( .IN1(\regf[24][11] ), .IN3(\regf[26][11] ), .IN2(
        \regf[25][11] ), .IN4(\regf[27][11] ), .S0(n1260), .S1(n1190), .Q(
        n2022) );
  MUX41X1 U2512 ( .IN1(\regf[20][11] ), .IN3(\regf[22][11] ), .IN2(
        \regf[21][11] ), .IN4(\regf[23][11] ), .S0(n1264), .S1(n1097), .Q(
        n2023) );
  MUX41X1 U2513 ( .IN1(\regf[16][11] ), .IN3(\regf[18][11] ), .IN2(
        \regf[17][11] ), .IN4(\regf[19][11] ), .S0(n1236), .S1(n1375), .Q(
        n2024) );
  MUX41X1 U2514 ( .IN1(\regf[12][11] ), .IN3(\regf[14][11] ), .IN2(
        \regf[13][11] ), .IN4(\regf[15][11] ), .S0(n1208), .S1(n1078), .Q(
        n2026) );
  MUX41X1 U2515 ( .IN1(\regf[8][11] ), .IN3(\regf[10][11] ), .IN2(
        \regf[9][11] ), .IN4(\regf[11][11] ), .S0(n1224), .S1(n1090), .Q(n2027) );
  MUX41X1 U2516 ( .IN1(\regf[4][11] ), .IN3(\regf[6][11] ), .IN2(\regf[5][11] ), .IN4(\regf[7][11] ), .S0(n1207), .S1(n1096), .Q(n2028) );
  MUX21X1 U2517 ( .IN1(n2030), .IN2(n2025), .S(n2381), .Q(rd_dataB[11]) );
  MUX41X1 U2518 ( .IN1(\regf[28][12] ), .IN3(\regf[30][12] ), .IN2(
        \regf[29][12] ), .IN4(\regf[31][12] ), .S0(n1265), .S1(n1139), .Q(
        n2031) );
  MUX41X1 U2519 ( .IN1(\regf[24][12] ), .IN3(\regf[26][12] ), .IN2(
        \regf[25][12] ), .IN4(\regf[27][12] ), .S0(n1208), .S1(n1112), .Q(
        n2032) );
  MUX41X1 U2520 ( .IN1(\regf[20][12] ), .IN3(\regf[22][12] ), .IN2(
        \regf[21][12] ), .IN4(\regf[23][12] ), .S0(n1265), .S1(n1137), .Q(
        n2033) );
  MUX41X1 U2521 ( .IN1(\regf[16][12] ), .IN3(\regf[18][12] ), .IN2(
        \regf[17][12] ), .IN4(\regf[19][12] ), .S0(n1265), .S1(n1156), .Q(
        n2034) );
  MUX41X1 U2522 ( .IN1(n2034), .IN3(n2032), .IN2(n2033), .IN4(n2031), .S0(
        n2376), .S1(n2370), .Q(n2035) );
  MUX41X1 U2523 ( .IN1(\regf[12][12] ), .IN3(\regf[14][12] ), .IN2(
        \regf[13][12] ), .IN4(\regf[15][12] ), .S0(n1258), .S1(n1133), .Q(
        n2036) );
  MUX41X1 U2524 ( .IN1(\regf[8][12] ), .IN3(\regf[10][12] ), .IN2(
        \regf[9][12] ), .IN4(\regf[11][12] ), .S0(n1225), .S1(n1375), .Q(n2037) );
  MUX41X1 U2525 ( .IN1(\regf[4][12] ), .IN3(\regf[6][12] ), .IN2(\regf[5][12] ), .IN4(\regf[7][12] ), .S0(n1208), .S1(n1181), .Q(n2038) );
  MUX41X1 U2526 ( .IN1(n2039), .IN3(n2037), .IN2(n2038), .IN4(n2036), .S0(
        n2376), .S1(n2370), .Q(n2040) );
  MUX21X1 U2527 ( .IN1(n2040), .IN2(n2035), .S(n2381), .Q(rd_dataB[12]) );
  MUX41X1 U2528 ( .IN1(\regf[28][13] ), .IN3(\regf[30][13] ), .IN2(
        \regf[29][13] ), .IN4(\regf[31][13] ), .S0(n1237), .S1(n1145), .Q(
        n2041) );
  MUX41X1 U2529 ( .IN1(\regf[24][13] ), .IN3(\regf[26][13] ), .IN2(
        \regf[25][13] ), .IN4(\regf[27][13] ), .S0(n1257), .S1(n1153), .Q(
        n2042) );
  MUX41X1 U2530 ( .IN1(\regf[20][13] ), .IN3(\regf[22][13] ), .IN2(
        \regf[21][13] ), .IN4(\regf[23][13] ), .S0(n1207), .S1(n1362), .Q(
        n2043) );
  MUX41X1 U2531 ( .IN1(\regf[16][13] ), .IN3(\regf[18][13] ), .IN2(
        \regf[17][13] ), .IN4(\regf[19][13] ), .S0(n1261), .S1(n1376), .Q(
        n2044) );
  MUX41X1 U2532 ( .IN1(n2044), .IN3(n2042), .IN2(n2043), .IN4(n2041), .S0(
        n2376), .S1(n2370), .Q(n2045) );
  MUX41X1 U2533 ( .IN1(\regf[12][13] ), .IN3(\regf[14][13] ), .IN2(
        \regf[13][13] ), .IN4(\regf[15][13] ), .S0(n1255), .S1(n1375), .Q(
        n2046) );
  MUX41X1 U2534 ( .IN1(\regf[8][13] ), .IN3(\regf[10][13] ), .IN2(
        \regf[9][13] ), .IN4(\regf[11][13] ), .S0(n1221), .S1(n1116), .Q(n2047) );
  MUX41X1 U2535 ( .IN1(\regf[4][13] ), .IN3(\regf[6][13] ), .IN2(\regf[5][13] ), .IN4(\regf[7][13] ), .S0(n1205), .S1(n1153), .Q(n2048) );
  MUX41X1 U2536 ( .IN1(\regf[28][14] ), .IN3(\regf[30][14] ), .IN2(
        \regf[29][14] ), .IN4(\regf[31][14] ), .S0(n1235), .S1(n1383), .Q(
        n2051) );
  MUX41X1 U2537 ( .IN1(\regf[24][14] ), .IN3(\regf[26][14] ), .IN2(
        \regf[25][14] ), .IN4(\regf[27][14] ), .S0(n1211), .S1(n1105), .Q(
        n2052) );
  MUX41X1 U2538 ( .IN1(\regf[20][14] ), .IN3(\regf[22][14] ), .IN2(
        \regf[21][14] ), .IN4(\regf[23][14] ), .S0(n1263), .S1(n1145), .Q(
        n2053) );
  MUX41X1 U2539 ( .IN1(\regf[16][14] ), .IN3(\regf[18][14] ), .IN2(
        \regf[17][14] ), .IN4(\regf[19][14] ), .S0(n1266), .S1(n1071), .Q(
        n2054) );
  MUX41X1 U2540 ( .IN1(\regf[12][14] ), .IN3(\regf[14][14] ), .IN2(
        \regf[13][14] ), .IN4(\regf[15][14] ), .S0(n1256), .S1(n1394), .Q(
        n2056) );
  MUX41X1 U2541 ( .IN1(\regf[8][14] ), .IN3(\regf[10][14] ), .IN2(
        \regf[9][14] ), .IN4(\regf[11][14] ), .S0(n1222), .S1(n1383), .Q(n2057) );
  MUX41X1 U2542 ( .IN1(\regf[4][14] ), .IN3(\regf[6][14] ), .IN2(\regf[5][14] ), .IN4(\regf[7][14] ), .S0(n1206), .S1(n1155), .Q(n2058) );
  MUX41X1 U2543 ( .IN1(n2059), .IN3(n2057), .IN2(n2058), .IN4(n2056), .S0(
        n2377), .S1(n2371), .Q(n2060) );
  MUX41X1 U2544 ( .IN1(\regf[28][15] ), .IN3(\regf[30][15] ), .IN2(
        \regf[29][15] ), .IN4(\regf[31][15] ), .S0(n1231), .S1(n1381), .Q(
        n2061) );
  MUX41X1 U2545 ( .IN1(\regf[24][15] ), .IN3(\regf[26][15] ), .IN2(
        \regf[25][15] ), .IN4(\regf[27][15] ), .S0(n1255), .S1(n1093), .Q(
        n2062) );
  MUX41X1 U2546 ( .IN1(\regf[20][15] ), .IN3(\regf[22][15] ), .IN2(
        \regf[21][15] ), .IN4(\regf[23][15] ), .S0(n1262), .S1(n1384), .Q(
        n2063) );
  MUX41X1 U2547 ( .IN1(\regf[16][15] ), .IN3(\regf[18][15] ), .IN2(
        \regf[17][15] ), .IN4(\regf[19][15] ), .S0(n1266), .S1(n1116), .Q(
        n2064) );
  MUX41X1 U2548 ( .IN1(\regf[12][15] ), .IN3(\regf[14][15] ), .IN2(
        \regf[13][15] ), .IN4(\regf[15][15] ), .S0(n1254), .S1(n1372), .Q(
        n2066) );
  MUX41X1 U2549 ( .IN1(\regf[8][15] ), .IN3(\regf[10][15] ), .IN2(
        \regf[9][15] ), .IN4(\regf[11][15] ), .S0(n1223), .S1(n1381), .Q(n2067) );
  MUX41X1 U2550 ( .IN1(\regf[4][15] ), .IN3(\regf[6][15] ), .IN2(\regf[5][15] ), .IN4(\regf[7][15] ), .S0(n1222), .S1(n1130), .Q(n2068) );
  MUX41X1 U2551 ( .IN1(\regf[28][16] ), .IN3(\regf[30][16] ), .IN2(
        \regf[29][16] ), .IN4(\regf[31][16] ), .S0(n1234), .S1(n1139), .Q(
        n2071) );
  MUX41X1 U2552 ( .IN1(\regf[24][16] ), .IN3(\regf[26][16] ), .IN2(
        \regf[25][16] ), .IN4(\regf[27][16] ), .S0(n1254), .S1(n1152), .Q(
        n2072) );
  MUX41X1 U2553 ( .IN1(\regf[20][16] ), .IN3(\regf[22][16] ), .IN2(
        \regf[21][16] ), .IN4(\regf[23][16] ), .S0(n1117), .S1(n1166), .Q(
        n2073) );
  MUX41X1 U2554 ( .IN1(\regf[16][16] ), .IN3(\regf[18][16] ), .IN2(
        \regf[17][16] ), .IN4(\regf[19][16] ), .S0(n1265), .S1(n1116), .Q(
        n2074) );
  MUX41X1 U2555 ( .IN1(n2074), .IN3(n2072), .IN2(n2073), .IN4(n2071), .S0(
        n2377), .S1(n2371), .Q(n2075) );
  MUX41X1 U2556 ( .IN1(\regf[12][16] ), .IN3(\regf[14][16] ), .IN2(
        \regf[13][16] ), .IN4(\regf[15][16] ), .S0(n1253), .S1(n1374), .Q(
        n2076) );
  MUX41X1 U2557 ( .IN1(\regf[8][16] ), .IN3(\regf[10][16] ), .IN2(
        \regf[9][16] ), .IN4(\regf[11][16] ), .S0(n1220), .S1(n1364), .Q(n2077) );
  MUX41X1 U2558 ( .IN1(\regf[4][16] ), .IN3(\regf[6][16] ), .IN2(\regf[5][16] ), .IN4(\regf[7][16] ), .S0(n1224), .S1(n1393), .Q(n2078) );
  MUX41X1 U2559 ( .IN1(n2079), .IN3(n2077), .IN2(n2078), .IN4(n2076), .S0(
        n2377), .S1(n2371), .Q(n2080) );
  MUX21X1 U2560 ( .IN1(n2080), .IN2(n2075), .S(n2381), .Q(rd_dataB[16]) );
  MUX41X1 U2561 ( .IN1(\regf[28][17] ), .IN3(\regf[30][17] ), .IN2(
        \regf[29][17] ), .IN4(\regf[31][17] ), .S0(n1232), .S1(n1363), .Q(
        n2081) );
  MUX41X1 U2562 ( .IN1(\regf[24][17] ), .IN3(\regf[26][17] ), .IN2(
        \regf[25][17] ), .IN4(\regf[27][17] ), .S0(n1256), .S1(n1109), .Q(
        n2082) );
  MUX41X1 U2563 ( .IN1(\regf[20][17] ), .IN3(\regf[22][17] ), .IN2(
        \regf[21][17] ), .IN4(\regf[23][17] ), .S0(n1268), .S1(n1393), .Q(
        n2083) );
  MUX41X1 U2564 ( .IN1(\regf[12][17] ), .IN3(\regf[14][17] ), .IN2(
        \regf[13][17] ), .IN4(\regf[15][17] ), .S0(n1211), .S1(n1154), .Q(
        n2086) );
  MUX41X1 U2565 ( .IN1(\regf[8][17] ), .IN3(\regf[10][17] ), .IN2(
        \regf[9][17] ), .IN4(\regf[11][17] ), .S0(n1236), .S1(n1375), .Q(n2087) );
  MUX41X1 U2566 ( .IN1(\regf[4][17] ), .IN3(\regf[6][17] ), .IN2(\regf[5][17] ), .IN4(\regf[7][17] ), .S0(n1223), .S1(n1355), .Q(n2088) );
  MUX41X1 U2567 ( .IN1(n2089), .IN3(n2087), .IN2(n2088), .IN4(n2086), .S0(
        n2377), .S1(n2371), .Q(n2090) );
  MUX41X1 U2568 ( .IN1(\regf[28][18] ), .IN3(\regf[30][18] ), .IN2(
        \regf[29][18] ), .IN4(\regf[31][18] ), .S0(n1254), .S1(n1396), .Q(
        n2091) );
  MUX41X1 U2569 ( .IN1(\regf[24][18] ), .IN3(\regf[26][18] ), .IN2(
        \regf[25][18] ), .IN4(\regf[27][18] ), .S0(n1250), .S1(n1390), .Q(
        n2092) );
  MUX41X1 U2570 ( .IN1(\regf[20][18] ), .IN3(\regf[22][18] ), .IN2(
        \regf[21][18] ), .IN4(\regf[23][18] ), .S0(n1273), .S1(n1133), .Q(
        n2093) );
  MUX41X1 U2571 ( .IN1(\regf[16][18] ), .IN3(\regf[18][18] ), .IN2(
        \regf[17][18] ), .IN4(\regf[19][18] ), .S0(n1252), .S1(n1392), .Q(
        n2094) );
  MUX41X1 U2572 ( .IN1(n2094), .IN3(n2092), .IN2(n2093), .IN4(n2091), .S0(
        n2377), .S1(n2371), .Q(n2095) );
  MUX41X1 U2573 ( .IN1(\regf[12][18] ), .IN3(\regf[14][18] ), .IN2(
        \regf[13][18] ), .IN4(\regf[15][18] ), .S0(n1262), .S1(n1374), .Q(
        n2096) );
  MUX41X1 U2574 ( .IN1(\regf[8][18] ), .IN3(\regf[10][18] ), .IN2(
        \regf[9][18] ), .IN4(\regf[11][18] ), .S0(n1265), .S1(n1372), .Q(n2097) );
  MUX41X1 U2575 ( .IN1(\regf[4][18] ), .IN3(\regf[6][18] ), .IN2(\regf[5][18] ), .IN4(\regf[7][18] ), .S0(n1227), .S1(n1396), .Q(n2098) );
  MUX41X1 U2576 ( .IN1(n2099), .IN3(n2097), .IN2(n2098), .IN4(n2096), .S0(
        n2377), .S1(n2371), .Q(n2100) );
  MUX41X1 U2577 ( .IN1(\regf[28][19] ), .IN3(\regf[30][19] ), .IN2(
        \regf[29][19] ), .IN4(\regf[31][19] ), .S0(n1249), .S1(n1391), .Q(
        n2101) );
  MUX41X1 U2578 ( .IN1(\regf[24][19] ), .IN3(\regf[26][19] ), .IN2(
        \regf[25][19] ), .IN4(\regf[27][19] ), .S0(n1117), .S1(n1391), .Q(
        n2102) );
  MUX41X1 U2579 ( .IN1(\regf[20][19] ), .IN3(\regf[22][19] ), .IN2(
        \regf[21][19] ), .IN4(\regf[23][19] ), .S0(n1274), .S1(n1105), .Q(
        n2103) );
  MUX41X1 U2580 ( .IN1(\regf[16][19] ), .IN3(\regf[18][19] ), .IN2(
        \regf[17][19] ), .IN4(\regf[19][19] ), .S0(n1206), .S1(n1090), .Q(
        n2104) );
  MUX41X1 U2581 ( .IN1(n2104), .IN3(n2102), .IN2(n2103), .IN4(n2101), .S0(
        n2377), .S1(n2371), .Q(n2105) );
  MUX41X1 U2582 ( .IN1(\regf[12][19] ), .IN3(\regf[14][19] ), .IN2(
        \regf[13][19] ), .IN4(\regf[15][19] ), .S0(n1274), .S1(n1354), .Q(
        n2106) );
  MUX41X1 U2583 ( .IN1(\regf[8][19] ), .IN3(\regf[10][19] ), .IN2(
        \regf[9][19] ), .IN4(\regf[11][19] ), .S0(n1230), .S1(n1354), .Q(n2107) );
  MUX41X1 U2584 ( .IN1(\regf[4][19] ), .IN3(\regf[6][19] ), .IN2(\regf[5][19] ), .IN4(\regf[7][19] ), .S0(n1267), .S1(n1372), .Q(n2108) );
  MUX41X1 U2585 ( .IN1(n2109), .IN3(n2107), .IN2(n2108), .IN4(n2106), .S0(
        n2377), .S1(n2371), .Q(n2110) );
  MUX41X1 U2586 ( .IN1(\regf[28][20] ), .IN3(\regf[30][20] ), .IN2(
        \regf[29][20] ), .IN4(\regf[31][20] ), .S0(n1207), .S1(n1140), .Q(
        n2111) );
  MUX41X1 U2587 ( .IN1(\regf[24][20] ), .IN3(\regf[26][20] ), .IN2(
        \regf[25][20] ), .IN4(\regf[27][20] ), .S0(n1210), .S1(n1375), .Q(
        n2112) );
  MUX41X1 U2588 ( .IN1(\regf[20][20] ), .IN3(\regf[22][20] ), .IN2(
        \regf[21][20] ), .IN4(\regf[23][20] ), .S0(n1246), .S1(n1109), .Q(
        n2113) );
  MUX41X1 U2589 ( .IN1(\regf[16][20] ), .IN3(\regf[18][20] ), .IN2(
        \regf[17][20] ), .IN4(\regf[19][20] ), .S0(n1207), .S1(n1137), .Q(
        n2114) );
  MUX41X1 U2590 ( .IN1(n2114), .IN3(n2112), .IN2(n2113), .IN4(n2111), .S0(
        n2378), .S1(n2372), .Q(n2115) );
  MUX41X1 U2591 ( .IN1(\regf[12][20] ), .IN3(\regf[14][20] ), .IN2(
        \regf[13][20] ), .IN4(\regf[15][20] ), .S0(n1206), .S1(n1140), .Q(
        n2116) );
  MUX41X1 U2592 ( .IN1(\regf[8][20] ), .IN3(\regf[10][20] ), .IN2(
        \regf[9][20] ), .IN4(\regf[11][20] ), .S0(n1231), .S1(n1355), .Q(n2117) );
  MUX41X1 U2593 ( .IN1(\regf[4][20] ), .IN3(\regf[6][20] ), .IN2(\regf[5][20] ), .IN4(\regf[7][20] ), .S0(n1208), .S1(n1381), .Q(n2118) );
  MUX41X1 U2594 ( .IN1(n2119), .IN3(n2117), .IN2(n2118), .IN4(n2116), .S0(
        n2378), .S1(n2372), .Q(n2120) );
  MUX21X1 U2595 ( .IN1(n2120), .IN2(n2115), .S(n2382), .Q(rd_dataB[20]) );
  MUX41X1 U2596 ( .IN1(\regf[28][21] ), .IN3(\regf[30][21] ), .IN2(
        \regf[29][21] ), .IN4(\regf[31][21] ), .S0(n1253), .S1(n1385), .Q(
        n2121) );
  MUX41X1 U2597 ( .IN1(\regf[24][21] ), .IN3(\regf[26][21] ), .IN2(
        \regf[25][21] ), .IN4(\regf[27][21] ), .S0(n1211), .S1(n1182), .Q(
        n2122) );
  MUX41X1 U2598 ( .IN1(\regf[20][21] ), .IN3(\regf[22][21] ), .IN2(
        \regf[21][21] ), .IN4(\regf[23][21] ), .S0(n1204), .S1(n1387), .Q(
        n2123) );
  MUX41X1 U2599 ( .IN1(\regf[16][21] ), .IN3(\regf[18][21] ), .IN2(
        \regf[17][21] ), .IN4(\regf[19][21] ), .S0(n1268), .S1(n1165), .Q(
        n2124) );
  MUX41X1 U2600 ( .IN1(\regf[12][21] ), .IN3(\regf[14][21] ), .IN2(
        \regf[13][21] ), .IN4(\regf[15][21] ), .S0(n1275), .S1(n1148), .Q(
        n2126) );
  MUX41X1 U2601 ( .IN1(\regf[8][21] ), .IN3(\regf[10][21] ), .IN2(
        \regf[9][21] ), .IN4(\regf[11][21] ), .S0(n1216), .S1(n1362), .Q(n2127) );
  MUX41X1 U2602 ( .IN1(\regf[4][21] ), .IN3(\regf[6][21] ), .IN2(\regf[5][21] ), .IN4(\regf[7][21] ), .S0(n1268), .S1(n1104), .Q(n2128) );
  MUX41X1 U2603 ( .IN1(n2129), .IN3(n2127), .IN2(n2128), .IN4(n2126), .S0(
        n2378), .S1(n2372), .Q(n2130) );
  MUX21X1 U2604 ( .IN1(n2130), .IN2(n2125), .S(n2382), .Q(rd_dataB[21]) );
  MUX41X1 U2605 ( .IN1(\regf[28][22] ), .IN3(\regf[30][22] ), .IN2(
        \regf[29][22] ), .IN4(\regf[31][22] ), .S0(n1209), .S1(n1170), .Q(
        n2131) );
  MUX41X1 U2606 ( .IN1(\regf[24][22] ), .IN3(\regf[26][22] ), .IN2(
        \regf[25][22] ), .IN4(\regf[27][22] ), .S0(n1212), .S1(n1381), .Q(
        n2132) );
  MUX41X1 U2607 ( .IN1(\regf[20][22] ), .IN3(\regf[22][22] ), .IN2(
        \regf[21][22] ), .IN4(\regf[23][22] ), .S0(n1211), .S1(n1143), .Q(
        n2133) );
  MUX41X1 U2608 ( .IN1(\regf[16][22] ), .IN3(\regf[18][22] ), .IN2(
        \regf[17][22] ), .IN4(\regf[19][22] ), .S0(n1269), .S1(n1148), .Q(
        n2134) );
  MUX41X1 U2609 ( .IN1(n2134), .IN3(n2132), .IN2(n2133), .IN4(n2131), .S0(
        n2378), .S1(n2372), .Q(n2135) );
  MUX41X1 U2610 ( .IN1(\regf[12][22] ), .IN3(\regf[14][22] ), .IN2(
        \regf[13][22] ), .IN4(\regf[15][22] ), .S0(n1209), .S1(n1366), .Q(
        n2136) );
  MUX41X1 U2611 ( .IN1(\regf[8][22] ), .IN3(\regf[10][22] ), .IN2(
        \regf[9][22] ), .IN4(\regf[11][22] ), .S0(n1265), .S1(n1157), .Q(n2137) );
  MUX41X1 U2612 ( .IN1(\regf[4][22] ), .IN3(\regf[6][22] ), .IN2(\regf[5][22] ), .IN4(\regf[7][22] ), .S0(n1269), .S1(n1358), .Q(n2138) );
  MUX41X1 U2613 ( .IN1(n2139), .IN3(n2137), .IN2(n2138), .IN4(n2136), .S0(
        n2378), .S1(n2372), .Q(n2140) );
  MUX21X1 U2614 ( .IN1(n2140), .IN2(n2135), .S(n2382), .Q(rd_dataB[22]) );
  MUX41X1 U2615 ( .IN1(\regf[28][23] ), .IN3(\regf[30][23] ), .IN2(
        \regf[29][23] ), .IN4(\regf[31][23] ), .S0(n1267), .S1(n1169), .Q(
        n2141) );
  MUX41X1 U2616 ( .IN1(\regf[20][23] ), .IN3(\regf[22][23] ), .IN2(
        \regf[21][23] ), .IN4(\regf[23][23] ), .S0(n1245), .S1(n1077), .Q(
        n2143) );
  MUX41X1 U2617 ( .IN1(\regf[16][23] ), .IN3(\regf[18][23] ), .IN2(
        \regf[17][23] ), .IN4(\regf[19][23] ), .S0(n1270), .S1(n1141), .Q(
        n2144) );
  MUX41X1 U2618 ( .IN1(n2144), .IN3(n2142), .IN2(n2143), .IN4(n2141), .S0(
        n2378), .S1(n2372), .Q(n2145) );
  MUX41X1 U2619 ( .IN1(\regf[12][23] ), .IN3(\regf[14][23] ), .IN2(
        \regf[13][23] ), .IN4(\regf[15][23] ), .S0(n1204), .S1(n1377), .Q(
        n2146) );
  MUX41X1 U2620 ( .IN1(\regf[8][23] ), .IN3(\regf[10][23] ), .IN2(
        \regf[9][23] ), .IN4(\regf[11][23] ), .S0(n1217), .S1(n1381), .Q(n2147) );
  MUX41X1 U2621 ( .IN1(\regf[4][23] ), .IN3(\regf[6][23] ), .IN2(\regf[5][23] ), .IN4(\regf[7][23] ), .S0(n1270), .S1(n1106), .Q(n2148) );
  MUX41X1 U2622 ( .IN1(n2149), .IN3(n2147), .IN2(n2148), .IN4(n2146), .S0(
        n2378), .S1(n2372), .Q(n2150) );
  MUX21X1 U2623 ( .IN1(n2150), .IN2(n2145), .S(n2382), .Q(rd_dataB[23]) );
  MUX41X1 U2624 ( .IN1(\regf[28][24] ), .IN3(\regf[30][24] ), .IN2(
        \regf[29][24] ), .IN4(\regf[31][24] ), .S0(n1266), .S1(n1167), .Q(
        n2151) );
  MUX41X1 U2625 ( .IN1(\regf[24][24] ), .IN3(\regf[26][24] ), .IN2(
        \regf[25][24] ), .IN4(\regf[27][24] ), .S0(n1214), .S1(n1145), .Q(
        n2152) );
  MUX41X1 U2626 ( .IN1(\regf[20][24] ), .IN3(\regf[22][24] ), .IN2(
        \regf[21][24] ), .IN4(\regf[23][24] ), .S0(n1125), .S1(n1164), .Q(
        n2153) );
  MUX41X1 U2627 ( .IN1(\regf[16][24] ), .IN3(\regf[18][24] ), .IN2(
        \regf[17][24] ), .IN4(\regf[19][24] ), .S0(n1271), .S1(n1384), .Q(
        n2154) );
  MUX41X1 U2628 ( .IN1(n2154), .IN3(n2152), .IN2(n2153), .IN4(n2151), .S0(
        n2378), .S1(n2372), .Q(n2155) );
  MUX41X1 U2629 ( .IN1(\regf[12][24] ), .IN3(\regf[14][24] ), .IN2(
        \regf[13][24] ), .IN4(\regf[15][24] ), .S0(n1205), .S1(n1392), .Q(
        n2156) );
  MUX41X1 U2630 ( .IN1(\regf[8][24] ), .IN3(\regf[10][24] ), .IN2(
        \regf[9][24] ), .IN4(\regf[11][24] ), .S0(n1232), .S1(n1107), .Q(n2157) );
  MUX41X1 U2631 ( .IN1(\regf[4][24] ), .IN3(\regf[6][24] ), .IN2(\regf[5][24] ), .IN4(\regf[7][24] ), .S0(n1271), .S1(n1190), .Q(n2158) );
  MUX41X1 U2632 ( .IN1(\regf[28][25] ), .IN3(\regf[30][25] ), .IN2(
        \regf[29][25] ), .IN4(\regf[31][25] ), .S0(n1205), .S1(n1092), .Q(
        n2161) );
  MUX41X1 U2633 ( .IN1(\regf[20][25] ), .IN3(\regf[22][25] ), .IN2(
        \regf[21][25] ), .IN4(\regf[23][25] ), .S0(n1275), .S1(n1171), .Q(
        n2163) );
  MUX41X1 U2634 ( .IN1(\regf[16][25] ), .IN3(\regf[18][25] ), .IN2(
        \regf[17][25] ), .IN4(\regf[19][25] ), .S0(n1272), .S1(n1088), .Q(
        n2164) );
  MUX41X1 U2635 ( .IN1(n2164), .IN3(n2162), .IN2(n2163), .IN4(n2161), .S0(
        n2378), .S1(n2372), .Q(n2165) );
  MUX41X1 U2636 ( .IN1(\regf[12][25] ), .IN3(\regf[14][25] ), .IN2(
        \regf[13][25] ), .IN4(\regf[15][25] ), .S0(n1207), .S1(n1142), .Q(
        n2166) );
  MUX41X1 U2637 ( .IN1(\regf[8][25] ), .IN3(\regf[10][25] ), .IN2(
        \regf[9][25] ), .IN4(\regf[11][25] ), .S0(n1233), .S1(n1156), .Q(n2167) );
  MUX41X1 U2638 ( .IN1(\regf[4][25] ), .IN3(\regf[6][25] ), .IN2(\regf[5][25] ), .IN4(\regf[7][25] ), .S0(n1272), .S1(n1390), .Q(n2168) );
  MUX41X1 U2639 ( .IN1(\regf[28][26] ), .IN3(\regf[30][26] ), .IN2(
        \regf[29][26] ), .IN4(\regf[31][26] ), .S0(n1267), .S1(n1142), .Q(
        n2171) );
  MUX41X1 U2640 ( .IN1(\regf[24][26] ), .IN3(\regf[26][26] ), .IN2(
        \regf[25][26] ), .IN4(\regf[27][26] ), .S0(n1216), .S1(n1384), .Q(
        n2172) );
  MUX41X1 U2641 ( .IN1(\regf[20][26] ), .IN3(\regf[22][26] ), .IN2(
        \regf[21][26] ), .IN4(\regf[23][26] ), .S0(n1205), .S1(n1167), .Q(
        n2173) );
  MUX41X1 U2642 ( .IN1(\regf[16][26] ), .IN3(\regf[18][26] ), .IN2(
        \regf[17][26] ), .IN4(\regf[19][26] ), .S0(n1273), .S1(n1097), .Q(
        n2174) );
  MUX41X1 U2643 ( .IN1(n2174), .IN3(n2172), .IN2(n2173), .IN4(n2171), .S0(
        n2379), .S1(n2373), .Q(n2175) );
  MUX41X1 U2644 ( .IN1(\regf[12][26] ), .IN3(\regf[14][26] ), .IN2(
        \regf[13][26] ), .IN4(\regf[15][26] ), .S0(n1208), .S1(n1110), .Q(
        n2176) );
  MUX41X1 U2645 ( .IN1(\regf[8][26] ), .IN3(\regf[10][26] ), .IN2(
        \regf[9][26] ), .IN4(\regf[11][26] ), .S0(n1234), .S1(n1089), .Q(n2177) );
  MUX41X1 U2646 ( .IN1(\regf[4][26] ), .IN3(\regf[6][26] ), .IN2(\regf[5][26] ), .IN4(\regf[7][26] ), .S0(n1273), .S1(n1191), .Q(n2178) );
  MUX21X1 U2647 ( .IN1(n2180), .IN2(n2175), .S(n2382), .Q(rd_dataB[26]) );
  MUX41X1 U2648 ( .IN1(\regf[28][27] ), .IN3(\regf[30][27] ), .IN2(
        \regf[29][27] ), .IN4(\regf[31][27] ), .S0(n1210), .S1(n1366), .Q(
        n2181) );
  MUX41X1 U2649 ( .IN1(\regf[24][27] ), .IN3(\regf[26][27] ), .IN2(
        \regf[25][27] ), .IN4(\regf[27][27] ), .S0(n1217), .S1(n1113), .Q(
        n2182) );
  MUX41X1 U2650 ( .IN1(\regf[20][27] ), .IN3(\regf[22][27] ), .IN2(
        \regf[21][27] ), .IN4(\regf[23][27] ), .S0(n1249), .S1(n1141), .Q(
        n2183) );
  MUX41X1 U2651 ( .IN1(\regf[16][27] ), .IN3(\regf[18][27] ), .IN2(
        \regf[17][27] ), .IN4(\regf[19][27] ), .S0(n1274), .S1(n1138), .Q(
        n2184) );
  MUX41X1 U2652 ( .IN1(n2184), .IN3(n2182), .IN2(n2183), .IN4(n2181), .S0(
        n2379), .S1(n2373), .Q(n2185) );
  MUX41X1 U2653 ( .IN1(\regf[12][27] ), .IN3(\regf[14][27] ), .IN2(
        \regf[13][27] ), .IN4(\regf[15][27] ), .S0(n1209), .S1(n1357), .Q(
        n2186) );
  MUX41X1 U2654 ( .IN1(\regf[8][27] ), .IN3(\regf[10][27] ), .IN2(
        \regf[9][27] ), .IN4(\regf[11][27] ), .S0(n1266), .S1(n1182), .Q(n2187) );
  MUX41X1 U2655 ( .IN1(\regf[4][27] ), .IN3(\regf[6][27] ), .IN2(\regf[5][27] ), .IN4(\regf[7][27] ), .S0(n1274), .S1(n1138), .Q(n2188) );
  MUX21X1 U2656 ( .IN1(n2190), .IN2(n2185), .S(n2382), .Q(rd_dataB[27]) );
  MUX41X1 U2657 ( .IN1(\regf[28][28] ), .IN3(\regf[30][28] ), .IN2(
        \regf[29][28] ), .IN4(\regf[31][28] ), .S0(n1211), .S1(n1143), .Q(
        n2191) );
  MUX41X1 U2658 ( .IN1(\regf[24][28] ), .IN3(\regf[26][28] ), .IN2(
        \regf[25][28] ), .IN4(\regf[27][28] ), .S0(n1218), .S1(n1393), .Q(
        n2192) );
  MUX41X1 U2659 ( .IN1(\regf[20][28] ), .IN3(\regf[22][28] ), .IN2(
        \regf[21][28] ), .IN4(\regf[23][28] ), .S0(n1252), .S1(n1358), .Q(
        n2193) );
  MUX41X1 U2660 ( .IN1(\regf[16][28] ), .IN3(\regf[18][28] ), .IN2(
        \regf[17][28] ), .IN4(\regf[19][28] ), .S0(n1275), .S1(n1107), .Q(
        n2194) );
  MUX41X1 U2661 ( .IN1(n2194), .IN3(n2192), .IN2(n2193), .IN4(n2191), .S0(
        n2379), .S1(n2373), .Q(n2195) );
  MUX41X1 U2662 ( .IN1(\regf[12][28] ), .IN3(\regf[14][28] ), .IN2(
        \regf[13][28] ), .IN4(\regf[15][28] ), .S0(n1210), .S1(n1363), .Q(
        n2196) );
  MUX41X1 U2663 ( .IN1(\regf[8][28] ), .IN3(\regf[10][28] ), .IN2(
        \regf[9][28] ), .IN4(\regf[11][28] ), .S0(n1235), .S1(n1385), .Q(n2197) );
  MUX41X1 U2664 ( .IN1(\regf[4][28] ), .IN3(\regf[6][28] ), .IN2(\regf[5][28] ), .IN4(\regf[7][28] ), .S0(n1275), .S1(n1116), .Q(n2198) );
  MUX41X1 U2665 ( .IN1(n2199), .IN3(n2197), .IN2(n2198), .IN4(n2196), .S0(
        n2379), .S1(n2373), .Q(n2200) );
  MUX41X1 U2666 ( .IN1(\regf[28][29] ), .IN3(\regf[30][29] ), .IN2(
        \regf[29][29] ), .IN4(\regf[31][29] ), .S0(n1268), .S1(n1171), .Q(
        n2201) );
  MUX41X1 U2667 ( .IN1(\regf[24][29] ), .IN3(\regf[26][29] ), .IN2(
        \regf[25][29] ), .IN4(\regf[27][29] ), .S0(n1219), .S1(n1163), .Q(
        n2202) );
  MUX41X1 U2668 ( .IN1(\regf[20][29] ), .IN3(\regf[22][29] ), .IN2(
        \regf[21][29] ), .IN4(\regf[23][29] ), .S0(n1251), .S1(n1095), .Q(
        n2203) );
  MUX41X1 U2669 ( .IN1(\regf[16][29] ), .IN3(\regf[18][29] ), .IN2(
        \regf[17][29] ), .IN4(\regf[19][29] ), .S0(n1210), .S1(n1077), .Q(
        n2204) );
  MUX41X1 U2670 ( .IN1(n2204), .IN3(n2202), .IN2(n2203), .IN4(n2201), .S0(
        n2379), .S1(n2373), .Q(n2205) );
  MUX41X1 U2671 ( .IN1(\regf[12][29] ), .IN3(\regf[14][29] ), .IN2(
        \regf[13][29] ), .IN4(\regf[15][29] ), .S0(n1211), .S1(n1396), .Q(
        n2206) );
  MUX41X1 U2672 ( .IN1(\regf[8][29] ), .IN3(\regf[10][29] ), .IN2(
        \regf[9][29] ), .IN4(\regf[11][29] ), .S0(n1204), .S1(n1165), .Q(n2207) );
  MUX41X1 U2673 ( .IN1(\regf[4][29] ), .IN3(\regf[6][29] ), .IN2(\regf[5][29] ), .IN4(\regf[7][29] ), .S0(n1206), .S1(n1359), .Q(n2208) );
  MUX41X1 U2674 ( .IN1(\regf[28][30] ), .IN3(\regf[30][30] ), .IN2(
        \regf[29][30] ), .IN4(\regf[31][30] ), .S0(n1211), .S1(n1382), .Q(
        n2211) );
  MUX41X1 U2675 ( .IN1(\regf[24][30] ), .IN3(\regf[26][30] ), .IN2(
        \regf[25][30] ), .IN4(\regf[27][30] ), .S0(n1204), .S1(n1113), .Q(
        n2212) );
  MUX41X1 U2676 ( .IN1(\regf[20][30] ), .IN3(\regf[22][30] ), .IN2(
        \regf[21][30] ), .IN4(\regf[23][30] ), .S0(n1269), .S1(n1391), .Q(
        n2213) );
  MUX41X1 U2677 ( .IN1(\regf[16][30] ), .IN3(\regf[18][30] ), .IN2(
        \regf[17][30] ), .IN4(\regf[19][30] ), .S0(n1263), .S1(n1188), .Q(
        n2214) );
  MUX41X1 U2678 ( .IN1(\regf[12][30] ), .IN3(\regf[14][30] ), .IN2(
        \regf[13][30] ), .IN4(\regf[15][30] ), .S0(n1269), .S1(n1188), .Q(
        n2216) );
  MUX41X1 U2679 ( .IN1(\regf[8][30] ), .IN3(\regf[10][30] ), .IN2(
        \regf[9][30] ), .IN4(\regf[11][30] ), .S0(n1212), .S1(n1374), .Q(n2217) );
  MUX41X1 U2680 ( .IN1(\regf[4][30] ), .IN3(\regf[6][30] ), .IN2(\regf[5][30] ), .IN4(\regf[7][30] ), .S0(n1117), .S1(n1094), .Q(n2218) );
  MUX41X1 U2681 ( .IN1(n2219), .IN3(n2217), .IN2(n2218), .IN4(n2216), .S0(
        n2379), .S1(n2373), .Q(n2220) );
  MUX41X1 U2682 ( .IN1(\regf[28][31] ), .IN3(\regf[30][31] ), .IN2(
        \regf[29][31] ), .IN4(\regf[31][31] ), .S0(n1204), .S1(n1384), .Q(
        n2221) );
  MUX41X1 U2683 ( .IN1(\regf[24][31] ), .IN3(\regf[26][31] ), .IN2(
        \regf[25][31] ), .IN4(\regf[27][31] ), .S0(n1205), .S1(n1137), .Q(
        n2222) );
  MUX41X1 U2684 ( .IN1(\regf[20][31] ), .IN3(\regf[22][31] ), .IN2(
        \regf[21][31] ), .IN4(\regf[23][31] ), .S0(n1208), .S1(n1364), .Q(
        n2223) );
  MUX41X1 U2685 ( .IN1(\regf[16][31] ), .IN3(\regf[18][31] ), .IN2(
        \regf[17][31] ), .IN4(\regf[19][31] ), .S0(n1265), .S1(n1387), .Q(
        n2224) );
  MUX41X1 U2686 ( .IN1(n2224), .IN3(n2222), .IN2(n2223), .IN4(n2221), .S0(
        n2379), .S1(n2373), .Q(n2225) );
  MUX41X1 U2687 ( .IN1(\regf[12][31] ), .IN3(\regf[14][31] ), .IN2(
        \regf[13][31] ), .IN4(\regf[15][31] ), .S0(n1270), .S1(n1130), .Q(
        n2226) );
  MUX41X1 U2688 ( .IN1(\regf[8][31] ), .IN3(\regf[10][31] ), .IN2(
        \regf[9][31] ), .IN4(\regf[11][31] ), .S0(n1213), .S1(n1137), .Q(n2227) );
  MUX41X1 U2689 ( .IN1(\regf[4][31] ), .IN3(\regf[6][31] ), .IN2(\regf[5][31] ), .IN4(\regf[7][31] ), .S0(n1265), .S1(n1163), .Q(n2228) );
  MUX41X1 U2690 ( .IN1(n2229), .IN3(n2227), .IN2(n2228), .IN4(n2226), .S0(
        n2379), .S1(n2373), .Q(n2230) );
  MUX21X1 U2691 ( .IN1(n2235), .IN2(n2236), .S(n1234), .Q(n2238) );
  NAND3X0 U2692 ( .IN1(\regf[3][30] ), .IN2(n1214), .IN3(n1189), .QN(n2237) );
  MUX21X1 U2693 ( .IN1(n2243), .IN2(n2244), .S(n1214), .Q(n2246) );
  MUX21X1 U2694 ( .IN1(n2247), .IN2(n2248), .S(n1235), .Q(n2250) );
  MUX21X1 U2695 ( .IN1(n2251), .IN2(n2252), .S(n1215), .Q(n2254) );
  NAND3X0 U2696 ( .IN1(\regf[3][25] ), .IN2(n1125), .IN3(n1187), .QN(n2257) );
  MUX21X1 U2697 ( .IN1(n2259), .IN2(n2260), .S(n1236), .Q(n2262) );
  MUX21X1 U2698 ( .IN1(n2263), .IN2(n2264), .S(n1217), .Q(n2266) );
  MUX21X1 U2699 ( .IN1(n2267), .IN2(n2268), .S(n1218), .Q(n2270) );
  MUX21X1 U2700 ( .IN1(n2271), .IN2(n2272), .S(n1237), .Q(n2274) );
  MUX21X1 U2701 ( .IN1(n2275), .IN2(n2276), .S(n1219), .Q(n2278) );
  MUX21X1 U2702 ( .IN1(n2279), .IN2(n2280), .S(n1231), .Q(n2282) );
  MUX21X1 U2703 ( .IN1(n2283), .IN2(n2284), .S(n1238), .Q(n2286) );
  MUX21X1 U2704 ( .IN1(n2287), .IN2(n2288), .S(n1237), .Q(n2290) );
  MUX21X1 U2705 ( .IN1(n2291), .IN2(n2292), .S(n1232), .Q(n2294) );
  NAND3X0 U2706 ( .IN1(\regf[3][16] ), .IN2(n1212), .IN3(n1392), .QN(n2293) );
  MUX21X1 U2707 ( .IN1(n2295), .IN2(n2296), .S(n1221), .Q(n2298) );
  NAND3X0 U2708 ( .IN1(\regf[3][15] ), .IN2(n1209), .IN3(n1189), .QN(n2297) );
  MUX21X1 U2709 ( .IN1(n2299), .IN2(n2300), .S(n1233), .Q(n2302) );
  NAND3X0 U2710 ( .IN1(\regf[3][13] ), .IN2(n1210), .IN3(n1186), .QN(n2305) );
  MUX21X1 U2711 ( .IN1(n2307), .IN2(n2308), .S(n1223), .Q(n2310) );
  NAND3X0 U2712 ( .IN1(\regf[3][10] ), .IN2(n1206), .IN3(n1187), .QN(n2317) );
  MUX21X1 U2713 ( .IN1(n2319), .IN2(n2320), .S(n1225), .Q(n2322) );
  MUX21X1 U2714 ( .IN1(n2323), .IN2(n2324), .S(n1220), .Q(n2326) );
  MUX21X1 U2715 ( .IN1(n2327), .IN2(n2328), .S(n1222), .Q(n2330) );
  NAND3X0 U2716 ( .IN1(\regf[3][6] ), .IN2(n1210), .IN3(n1364), .QN(n2333) );
  MUX21X1 U2717 ( .IN1(n2339), .IN2(n2340), .S(n1226), .Q(n2342) );
  MUX21X1 U2718 ( .IN1(n2351), .IN2(n2352), .S(n1235), .Q(n2354) );
  NAND3X0 U2719 ( .IN1(\regf[3][1] ), .IN2(n1216), .IN3(n1186), .QN(n2353) );
  MUX21X1 U2720 ( .IN1(n2355), .IN2(n2356), .S(n1230), .Q(n2358) );
  INVX0 U2721 ( .INP(N16), .ZN(n2359) );
  INVX0 U2722 ( .INP(N16), .ZN(n2360) );
  DELLN1X2 U2723 ( .INP(N17), .Z(n2367) );
  DELLN1X2 U2724 ( .INP(N18), .Z(n2369) );
  DELLN1X2 U2725 ( .INP(N18), .Z(n2370) );
  DELLN1X2 U2726 ( .INP(N18), .Z(n2371) );
  DELLN1X2 U2727 ( .INP(N18), .Z(n2372) );
  DELLN1X2 U2728 ( .INP(N18), .Z(n2373) );
  DELLN1X2 U2729 ( .INP(N20), .Z(n2382) );
  DELLN1X2 U2730 ( .INP(N19), .Z(n2379) );
  NAND2X0 U2731 ( .IN1(n71), .IN2(n51), .QN(n78) );
  NAND2X0 U2732 ( .IN1(n71), .IN2(n49), .QN(n77) );
  NAND2X0 U2733 ( .IN1(n71), .IN2(n47), .QN(n76) );
  NAND2X0 U2734 ( .IN1(n71), .IN2(n45), .QN(n75) );
  NAND2X0 U2735 ( .IN1(n71), .IN2(n36), .QN(n70) );
  INVX0 U2736 ( .INP(n74), .ZN(n2402) );
  NAND2X0 U2737 ( .IN1(n71), .IN2(n43), .QN(n74) );
  NAND2X0 U2738 ( .IN1(n53), .IN2(n49), .QN(n59) );
  NAND2X0 U2739 ( .IN1(n53), .IN2(n47), .QN(n58) );
  NAND2X0 U2740 ( .IN1(n53), .IN2(n45), .QN(n57) );
  NAND2X0 U2741 ( .IN1(n53), .IN2(n51), .QN(n60) );
  INVX0 U2742 ( .INP(n73), .ZN(n2407) );
  NAND2X0 U2743 ( .IN1(n71), .IN2(n41), .QN(n73) );
  INVX0 U2744 ( .INP(n72), .ZN(n2412) );
  NAND2X0 U2745 ( .IN1(n71), .IN2(n38), .QN(n72) );
  INVX0 U2746 ( .INP(n56), .ZN(n2477) );
  NAND2X0 U2747 ( .IN1(n53), .IN2(n2383), .QN(n56) );
  NAND2X0 U2748 ( .IN1(n53), .IN2(n36), .QN(n52) );
  INVX0 U2749 ( .INP(n55), .ZN(n2482) );
  NAND2X0 U2750 ( .IN1(n53), .IN2(n41), .QN(n55) );
  INVX0 U2751 ( .INP(n54), .ZN(n2487) );
  NAND2X0 U2752 ( .IN1(n53), .IN2(n38), .QN(n54) );
  NAND2X0 U2753 ( .IN1(n49), .IN2(n39), .QN(n48) );
  NAND2X0 U2754 ( .IN1(n47), .IN2(n39), .QN(n46) );
  NAND2X0 U2755 ( .IN1(n45), .IN2(n39), .QN(n44) );
  NAND2X0 U2756 ( .IN1(n51), .IN2(n39), .QN(n50) );
  INVX0 U2757 ( .INP(n42), .ZN(n2512) );
  NAND2X0 U2758 ( .IN1(n2383), .IN2(n39), .QN(n42) );
  INVX0 U2759 ( .INP(n37), .ZN(n2522) );
  NAND2X0 U2760 ( .IN1(n38), .IN2(n39), .QN(n37) );
  INVX0 U2761 ( .INP(n40), .ZN(n2517) );
  NAND2X0 U2762 ( .IN1(n41), .IN2(n39), .QN(n40) );
  INVX0 U2763 ( .INP(wr_addr[4]), .ZN(n2711) );
  NAND2X0 U2764 ( .IN1(n62), .IN2(n36), .QN(n61) );
  NAND2X0 U2765 ( .IN1(n62), .IN2(n38), .QN(n63) );
  NAND2X0 U2766 ( .IN1(n62), .IN2(n41), .QN(n64) );
  NAND2X0 U2767 ( .IN1(n62), .IN2(n43), .QN(n65) );
  NAND2X0 U2768 ( .IN1(n62), .IN2(n45), .QN(n66) );
  NAND2X0 U2769 ( .IN1(n62), .IN2(n47), .QN(n67) );
  NAND2X0 U2770 ( .IN1(n62), .IN2(n49), .QN(n68) );
  NOR3X0 U2771 ( .IN1(n2714), .IN2(wr_addr[2]), .IN3(n2713), .QN(n2383) );
  INVX0 U2772 ( .INP(wr_addr[1]), .ZN(n2713) );
  INVX0 U2773 ( .INP(wr_addr[0]), .ZN(n2714) );
  INVX0 U2774 ( .INP(n2386), .ZN(n2384) );
  INVX0 U2775 ( .INP(n2387), .ZN(n2385) );
  INVX0 U2776 ( .INP(n2390), .ZN(n2388) );
  INVX0 U2777 ( .INP(n2391), .ZN(n2389) );
  INVX0 U2778 ( .INP(n2394), .ZN(n2392) );
  INVX0 U2779 ( .INP(n2395), .ZN(n2393) );
  INVX0 U2780 ( .INP(n2398), .ZN(n2396) );
  INVX0 U2781 ( .INP(n2399), .ZN(n2397) );
  INVX0 U2782 ( .INP(n2402), .ZN(n2400) );
  INVX0 U2783 ( .INP(n2402), .ZN(n2401) );
  INVX0 U2784 ( .INP(n2407), .ZN(n2405) );
  INVX0 U2785 ( .INP(n2407), .ZN(n2406) );
  INVX0 U2786 ( .INP(n2412), .ZN(n2410) );
  INVX0 U2787 ( .INP(n2412), .ZN(n2411) );
  INVX0 U2788 ( .INP(n2417), .ZN(n2415) );
  INVX0 U2789 ( .INP(n2418), .ZN(n2416) );
  INVX0 U2790 ( .INP(n2421), .ZN(n2419) );
  INVX0 U2791 ( .INP(n2421), .ZN(n2420) );
  INVX0 U2792 ( .INP(n2426), .ZN(n2424) );
  INVX0 U2793 ( .INP(n2426), .ZN(n2425) );
  INVX0 U2794 ( .INP(n2431), .ZN(n2429) );
  INVX0 U2795 ( .INP(n2431), .ZN(n2430) );
  INVX0 U2796 ( .INP(n2436), .ZN(n2434) );
  INVX0 U2797 ( .INP(n2436), .ZN(n2435) );
  INVX0 U2798 ( .INP(n2441), .ZN(n2439) );
  INVX0 U2799 ( .INP(n2441), .ZN(n2440) );
  INVX0 U2800 ( .INP(n2446), .ZN(n2444) );
  INVX0 U2801 ( .INP(n2446), .ZN(n2445) );
  INVX0 U2802 ( .INP(n2451), .ZN(n2449) );
  INVX0 U2803 ( .INP(n2451), .ZN(n2450) );
  INVX0 U2804 ( .INP(n2456), .ZN(n2454) );
  INVX0 U2805 ( .INP(n2456), .ZN(n2455) );
  INVX0 U2806 ( .INP(n2461), .ZN(n2459) );
  INVX0 U2807 ( .INP(n2462), .ZN(n2460) );
  INVX0 U2808 ( .INP(n2465), .ZN(n2463) );
  INVX0 U2809 ( .INP(n2466), .ZN(n2464) );
  INVX0 U2810 ( .INP(n2469), .ZN(n2467) );
  INVX0 U2811 ( .INP(n2470), .ZN(n2468) );
  INVX0 U2812 ( .INP(n2473), .ZN(n2471) );
  INVX0 U2813 ( .INP(n2474), .ZN(n2472) );
  INVX0 U2814 ( .INP(n2477), .ZN(n2475) );
  INVX0 U2815 ( .INP(n2477), .ZN(n2476) );
  INVX0 U2816 ( .INP(n2482), .ZN(n2480) );
  INVX0 U2817 ( .INP(n2482), .ZN(n2481) );
  INVX0 U2818 ( .INP(n2487), .ZN(n2485) );
  INVX0 U2819 ( .INP(n2487), .ZN(n2486) );
  INVX0 U2820 ( .INP(n2492), .ZN(n2490) );
  INVX0 U2821 ( .INP(n2493), .ZN(n2491) );
  INVX0 U2822 ( .INP(n2496), .ZN(n2494) );
  INVX0 U2823 ( .INP(n2497), .ZN(n2495) );
  INVX0 U2824 ( .INP(n2500), .ZN(n2498) );
  INVX0 U2825 ( .INP(n2501), .ZN(n2499) );
  INVX0 U2826 ( .INP(n2504), .ZN(n2502) );
  INVX0 U2827 ( .INP(n2505), .ZN(n2503) );
  INVX0 U2828 ( .INP(n2508), .ZN(n2506) );
  INVX0 U2829 ( .INP(n2509), .ZN(n2507) );
  INVX0 U2830 ( .INP(n2512), .ZN(n2510) );
  INVX0 U2831 ( .INP(n2512), .ZN(n2511) );
  INVX0 U2832 ( .INP(n2517), .ZN(n2515) );
  INVX0 U2833 ( .INP(n2517), .ZN(n2516) );
  INVX0 U2834 ( .INP(n2522), .ZN(n2520) );
  INVX0 U2835 ( .INP(n2522), .ZN(n2521) );
endmodule

