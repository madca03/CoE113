`timescale 1ns/1ps
module rf ( clk, rst_n, rd_addrA, rd_addrB, rd_dataA, rd_dataB, wr_en, wr_addr, 
        wr_data );
  input [4:0] rd_addrA;
  input [4:0] rd_addrB;
  output [31:0] rd_dataA;
  output [31:0] rd_dataB;
  input [4:0] wr_addr;
  input [31:0] wr_data;
  input clk, rst_n, wr_en;
  wire   N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393;
  wire   [31:0] reg2;
  wire   [31:0] reg3;
  wire   [31:0] reg4;
  wire   [31:0] reg5;
  wire   [31:0] reg6;
  wire   [31:0] reg7;
  wire   [31:0] reg8;
  wire   [31:0] reg9;
  wire   [31:0] reg10;
  wire   [31:0] reg11;
  wire   [31:0] reg12;
  wire   [31:0] reg13;
  wire   [31:0] reg14;
  wire   [31:0] reg15;
  wire   [31:0] reg16;
  wire   [31:0] reg17;
  wire   [31:0] reg18;
  wire   [31:0] reg19;
  wire   [31:0] reg20;
  wire   [31:0] reg21;
  wire   [31:0] reg22;
  wire   [31:0] reg23;
  wire   [31:0] reg24;
  wire   [31:0] reg25;
  wire   [31:0] reg26;
  wire   [31:0] reg27;
  wire   [31:0] reg28;
  wire   [31:0] reg29;
  wire   [31:0] reg30;
  wire   [31:0] reg31;
  wire   [31:0] reg32;
  assign N11 = rd_addrA[0];
  assign N12 = rd_addrA[1];
  assign N13 = rd_addrA[2];
  assign N14 = rd_addrA[3];
  assign N15 = rd_addrA[4];
  assign N16 = rd_addrB[0];
  assign N17 = rd_addrB[1];
  assign N18 = rd_addrB[2];
  assign N19 = rd_addrB[3];
  assign N20 = rd_addrB[4];

  DFFARX1 \regf_reg[31][31]  ( .D(n1070), .CLK(clk), .RSTB(n2382), .Q(
        reg32[31]) );
  DFFARX1 \regf_reg[31][30]  ( .D(n1069), .CLK(clk), .RSTB(n2382), .Q(
        reg32[30]) );
  DFFARX1 \regf_reg[31][29]  ( .D(n1068), .CLK(clk), .RSTB(n2382), .Q(
        reg32[29]) );
  DFFARX1 \regf_reg[31][28]  ( .D(n1067), .CLK(clk), .RSTB(n2382), .Q(
        reg32[28]) );
  DFFARX1 \regf_reg[31][27]  ( .D(n1066), .CLK(clk), .RSTB(n2382), .Q(
        reg32[27]) );
  DFFARX1 \regf_reg[31][26]  ( .D(n1065), .CLK(clk), .RSTB(n2382), .Q(
        reg32[26]) );
  DFFARX1 \regf_reg[31][25]  ( .D(n1064), .CLK(clk), .RSTB(n2382), .Q(
        reg32[25]) );
  DFFARX1 \regf_reg[31][24]  ( .D(n1063), .CLK(clk), .RSTB(n2382), .Q(
        reg32[24]) );
  DFFARX1 \regf_reg[31][23]  ( .D(n1062), .CLK(clk), .RSTB(n2381), .Q(
        reg32[23]) );
  DFFARX1 \regf_reg[31][22]  ( .D(n1061), .CLK(clk), .RSTB(n2381), .Q(
        reg32[22]) );
  DFFARX1 \regf_reg[31][21]  ( .D(n1060), .CLK(clk), .RSTB(n2381), .Q(
        reg32[21]) );
  DFFARX1 \regf_reg[31][20]  ( .D(n1059), .CLK(clk), .RSTB(n2381), .Q(
        reg32[20]) );
  DFFARX1 \regf_reg[31][19]  ( .D(n1058), .CLK(clk), .RSTB(n2381), .Q(
        reg32[19]) );
  DFFARX1 \regf_reg[31][18]  ( .D(n1057), .CLK(clk), .RSTB(n2381), .Q(
        reg32[18]) );
  DFFARX1 \regf_reg[31][17]  ( .D(n1056), .CLK(clk), .RSTB(n2381), .Q(
        reg32[17]) );
  DFFARX1 \regf_reg[31][16]  ( .D(n1055), .CLK(clk), .RSTB(n2381), .Q(
        reg32[16]) );
  DFFARX1 \regf_reg[31][15]  ( .D(n1054), .CLK(clk), .RSTB(n2381), .Q(
        reg32[15]) );
  DFFARX1 \regf_reg[31][14]  ( .D(n1053), .CLK(clk), .RSTB(n2381), .Q(
        reg32[14]) );
  DFFARX1 \regf_reg[31][13]  ( .D(n1052), .CLK(clk), .RSTB(n2381), .Q(
        reg32[13]) );
  DFFARX1 \regf_reg[31][12]  ( .D(n1051), .CLK(clk), .RSTB(n2381), .Q(
        reg32[12]) );
  DFFARX1 \regf_reg[31][11]  ( .D(n1050), .CLK(clk), .RSTB(n2380), .Q(
        reg32[11]) );
  DFFARX1 \regf_reg[31][10]  ( .D(n1049), .CLK(clk), .RSTB(n2380), .Q(
        reg32[10]) );
  DFFARX1 \regf_reg[31][9]  ( .D(n1048), .CLK(clk), .RSTB(n2380), .Q(reg32[9])
         );
  DFFARX1 \regf_reg[31][8]  ( .D(n1047), .CLK(clk), .RSTB(n2380), .Q(reg32[8])
         );
  DFFARX1 \regf_reg[31][7]  ( .D(n1046), .CLK(clk), .RSTB(n2380), .Q(reg32[7])
         );
  DFFARX1 \regf_reg[31][6]  ( .D(n1045), .CLK(clk), .RSTB(n2380), .Q(reg32[6])
         );
  DFFARX1 \regf_reg[31][5]  ( .D(n1044), .CLK(clk), .RSTB(n2380), .Q(reg32[5])
         );
  DFFARX1 \regf_reg[31][4]  ( .D(n1043), .CLK(clk), .RSTB(n2380), .Q(reg32[4])
         );
  DFFARX1 \regf_reg[31][3]  ( .D(n1042), .CLK(clk), .RSTB(n2380), .Q(reg32[3])
         );
  DFFARX1 \regf_reg[31][2]  ( .D(n1041), .CLK(clk), .RSTB(n2380), .Q(reg32[2])
         );
  DFFARX1 \regf_reg[31][1]  ( .D(n1040), .CLK(clk), .RSTB(n2380), .Q(reg32[1])
         );
  DFFARX1 \regf_reg[31][0]  ( .D(n1039), .CLK(clk), .RSTB(n2380), .Q(reg32[0])
         );
  DFFARX1 \regf_reg[30][31]  ( .D(n1038), .CLK(clk), .RSTB(n2379), .Q(
        reg31[31]) );
  DFFARX1 \regf_reg[30][30]  ( .D(n1037), .CLK(clk), .RSTB(n2379), .Q(
        reg31[30]) );
  DFFARX1 \regf_reg[30][29]  ( .D(n1036), .CLK(clk), .RSTB(n2379), .Q(
        reg31[29]) );
  DFFARX1 \regf_reg[30][28]  ( .D(n1035), .CLK(clk), .RSTB(n2379), .Q(
        reg31[28]) );
  DFFARX1 \regf_reg[30][27]  ( .D(n1034), .CLK(clk), .RSTB(n2379), .Q(
        reg31[27]) );
  DFFARX1 \regf_reg[30][26]  ( .D(n1033), .CLK(clk), .RSTB(n2379), .Q(
        reg31[26]) );
  DFFARX1 \regf_reg[30][25]  ( .D(n1032), .CLK(clk), .RSTB(n2379), .Q(
        reg31[25]) );
  DFFARX1 \regf_reg[30][24]  ( .D(n1031), .CLK(clk), .RSTB(n2379), .Q(
        reg31[24]) );
  DFFARX1 \regf_reg[30][23]  ( .D(n1030), .CLK(clk), .RSTB(n2379), .Q(
        reg31[23]) );
  DFFARX1 \regf_reg[30][22]  ( .D(n1029), .CLK(clk), .RSTB(n2379), .Q(
        reg31[22]) );
  DFFARX1 \regf_reg[30][21]  ( .D(n1028), .CLK(clk), .RSTB(n2379), .Q(
        reg31[21]) );
  DFFARX1 \regf_reg[30][20]  ( .D(n1027), .CLK(clk), .RSTB(n2379), .Q(
        reg31[20]) );
  DFFARX1 \regf_reg[30][19]  ( .D(n1026), .CLK(clk), .RSTB(n2378), .Q(
        reg31[19]) );
  DFFARX1 \regf_reg[30][18]  ( .D(n1025), .CLK(clk), .RSTB(n2378), .Q(
        reg31[18]) );
  DFFARX1 \regf_reg[30][17]  ( .D(n1024), .CLK(clk), .RSTB(n2378), .Q(
        reg31[17]) );
  DFFARX1 \regf_reg[30][16]  ( .D(n1023), .CLK(clk), .RSTB(n2378), .Q(
        reg31[16]) );
  DFFARX1 \regf_reg[30][15]  ( .D(n1022), .CLK(clk), .RSTB(n2378), .Q(
        reg31[15]) );
  DFFARX1 \regf_reg[30][14]  ( .D(n1021), .CLK(clk), .RSTB(n2378), .Q(
        reg31[14]) );
  DFFARX1 \regf_reg[30][13]  ( .D(n1020), .CLK(clk), .RSTB(n2378), .Q(
        reg31[13]) );
  DFFARX1 \regf_reg[30][12]  ( .D(n1019), .CLK(clk), .RSTB(n2378), .Q(
        reg31[12]) );
  DFFARX1 \regf_reg[30][11]  ( .D(n1018), .CLK(clk), .RSTB(n2378), .Q(
        reg31[11]) );
  DFFARX1 \regf_reg[30][10]  ( .D(n1017), .CLK(clk), .RSTB(n2378), .Q(
        reg31[10]) );
  DFFARX1 \regf_reg[30][9]  ( .D(n1016), .CLK(clk), .RSTB(n2378), .Q(reg31[9])
         );
  DFFARX1 \regf_reg[30][8]  ( .D(n1015), .CLK(clk), .RSTB(n2378), .Q(reg31[8])
         );
  DFFARX1 \regf_reg[30][7]  ( .D(n1014), .CLK(clk), .RSTB(n2377), .Q(reg31[7])
         );
  DFFARX1 \regf_reg[30][6]  ( .D(n1013), .CLK(clk), .RSTB(n2377), .Q(reg31[6])
         );
  DFFARX1 \regf_reg[30][5]  ( .D(n1012), .CLK(clk), .RSTB(n2377), .Q(reg31[5])
         );
  DFFARX1 \regf_reg[30][4]  ( .D(n1011), .CLK(clk), .RSTB(n2377), .Q(reg31[4])
         );
  DFFARX1 \regf_reg[30][3]  ( .D(n1010), .CLK(clk), .RSTB(n2377), .Q(reg31[3])
         );
  DFFARX1 \regf_reg[30][2]  ( .D(n1009), .CLK(clk), .RSTB(n2377), .Q(reg31[2])
         );
  DFFARX1 \regf_reg[30][1]  ( .D(n1008), .CLK(clk), .RSTB(n2377), .Q(reg31[1])
         );
  DFFARX1 \regf_reg[30][0]  ( .D(n1007), .CLK(clk), .RSTB(n2377), .Q(reg31[0])
         );
  DFFARX1 \regf_reg[29][31]  ( .D(n1006), .CLK(clk), .RSTB(n2377), .Q(
        reg30[31]) );
  DFFARX1 \regf_reg[29][30]  ( .D(n1005), .CLK(clk), .RSTB(n2377), .Q(
        reg30[30]) );
  DFFARX1 \regf_reg[29][29]  ( .D(n1004), .CLK(clk), .RSTB(n2377), .Q(
        reg30[29]) );
  DFFARX1 \regf_reg[29][28]  ( .D(n1003), .CLK(clk), .RSTB(n2377), .Q(
        reg30[28]) );
  DFFARX1 \regf_reg[29][27]  ( .D(n1002), .CLK(clk), .RSTB(n2376), .Q(
        reg30[27]) );
  DFFARX1 \regf_reg[29][26]  ( .D(n1001), .CLK(clk), .RSTB(n2376), .Q(
        reg30[26]) );
  DFFARX1 \regf_reg[29][25]  ( .D(n1000), .CLK(clk), .RSTB(n2376), .Q(
        reg30[25]) );
  DFFARX1 \regf_reg[29][24]  ( .D(n999), .CLK(clk), .RSTB(n2376), .Q(reg30[24]) );
  DFFARX1 \regf_reg[29][23]  ( .D(n998), .CLK(clk), .RSTB(n2376), .Q(reg30[23]) );
  DFFARX1 \regf_reg[29][22]  ( .D(n997), .CLK(clk), .RSTB(n2376), .Q(reg30[22]) );
  DFFARX1 \regf_reg[29][21]  ( .D(n996), .CLK(clk), .RSTB(n2376), .Q(reg30[21]) );
  DFFARX1 \regf_reg[29][20]  ( .D(n995), .CLK(clk), .RSTB(n2376), .Q(reg30[20]) );
  DFFARX1 \regf_reg[29][19]  ( .D(n994), .CLK(clk), .RSTB(n2376), .Q(reg30[19]) );
  DFFARX1 \regf_reg[29][18]  ( .D(n993), .CLK(clk), .RSTB(n2376), .Q(reg30[18]) );
  DFFARX1 \regf_reg[29][17]  ( .D(n992), .CLK(clk), .RSTB(n2376), .Q(reg30[17]) );
  DFFARX1 \regf_reg[29][16]  ( .D(n991), .CLK(clk), .RSTB(n2376), .Q(reg30[16]) );
  DFFARX1 \regf_reg[29][15]  ( .D(n990), .CLK(clk), .RSTB(n2375), .Q(reg30[15]) );
  DFFARX1 \regf_reg[29][14]  ( .D(n989), .CLK(clk), .RSTB(n2375), .Q(reg30[14]) );
  DFFARX1 \regf_reg[29][13]  ( .D(n988), .CLK(clk), .RSTB(n2375), .Q(reg30[13]) );
  DFFARX1 \regf_reg[29][12]  ( .D(n987), .CLK(clk), .RSTB(n2375), .Q(reg30[12]) );
  DFFARX1 \regf_reg[29][11]  ( .D(n986), .CLK(clk), .RSTB(n2375), .Q(reg30[11]) );
  DFFARX1 \regf_reg[29][10]  ( .D(n985), .CLK(clk), .RSTB(n2375), .Q(reg30[10]) );
  DFFARX1 \regf_reg[29][9]  ( .D(n984), .CLK(clk), .RSTB(n2375), .Q(reg30[9])
         );
  DFFARX1 \regf_reg[29][8]  ( .D(n983), .CLK(clk), .RSTB(n2375), .Q(reg30[8])
         );
  DFFARX1 \regf_reg[29][7]  ( .D(n982), .CLK(clk), .RSTB(n2375), .Q(reg30[7])
         );
  DFFARX1 \regf_reg[29][6]  ( .D(n981), .CLK(clk), .RSTB(n2375), .Q(reg30[6])
         );
  DFFARX1 \regf_reg[29][5]  ( .D(n980), .CLK(clk), .RSTB(n2375), .Q(reg30[5])
         );
  DFFARX1 \regf_reg[29][4]  ( .D(n979), .CLK(clk), .RSTB(n2375), .Q(reg30[4])
         );
  DFFARX1 \regf_reg[29][3]  ( .D(n978), .CLK(clk), .RSTB(n2374), .Q(reg30[3])
         );
  DFFARX1 \regf_reg[29][2]  ( .D(n977), .CLK(clk), .RSTB(n2374), .Q(reg30[2])
         );
  DFFARX1 \regf_reg[29][1]  ( .D(n976), .CLK(clk), .RSTB(n2374), .Q(reg30[1])
         );
  DFFARX1 \regf_reg[29][0]  ( .D(n975), .CLK(clk), .RSTB(n2374), .Q(reg30[0])
         );
  DFFARX1 \regf_reg[28][31]  ( .D(n974), .CLK(clk), .RSTB(n2374), .Q(reg29[31]) );
  DFFARX1 \regf_reg[28][30]  ( .D(n973), .CLK(clk), .RSTB(n2374), .Q(reg29[30]) );
  DFFARX1 \regf_reg[28][29]  ( .D(n972), .CLK(clk), .RSTB(n2374), .Q(reg29[29]) );
  DFFARX1 \regf_reg[28][28]  ( .D(n971), .CLK(clk), .RSTB(n2374), .Q(reg29[28]) );
  DFFARX1 \regf_reg[28][27]  ( .D(n970), .CLK(clk), .RSTB(n2374), .Q(reg29[27]) );
  DFFARX1 \regf_reg[28][26]  ( .D(n969), .CLK(clk), .RSTB(n2374), .Q(reg29[26]) );
  DFFARX1 \regf_reg[28][25]  ( .D(n968), .CLK(clk), .RSTB(n2374), .Q(reg29[25]) );
  DFFARX1 \regf_reg[28][24]  ( .D(n967), .CLK(clk), .RSTB(n2374), .Q(reg29[24]) );
  DFFARX1 \regf_reg[28][23]  ( .D(n966), .CLK(clk), .RSTB(n2373), .Q(reg29[23]) );
  DFFARX1 \regf_reg[28][22]  ( .D(n965), .CLK(clk), .RSTB(n2373), .Q(reg29[22]) );
  DFFARX1 \regf_reg[28][21]  ( .D(n964), .CLK(clk), .RSTB(n2373), .Q(reg29[21]) );
  DFFARX1 \regf_reg[28][20]  ( .D(n963), .CLK(clk), .RSTB(n2373), .Q(reg29[20]) );
  DFFARX1 \regf_reg[28][19]  ( .D(n962), .CLK(clk), .RSTB(n2373), .Q(reg29[19]) );
  DFFARX1 \regf_reg[28][18]  ( .D(n961), .CLK(clk), .RSTB(n2373), .Q(reg29[18]) );
  DFFARX1 \regf_reg[28][17]  ( .D(n960), .CLK(clk), .RSTB(n2373), .Q(reg29[17]) );
  DFFARX1 \regf_reg[28][16]  ( .D(n959), .CLK(clk), .RSTB(n2373), .Q(reg29[16]) );
  DFFARX1 \regf_reg[28][15]  ( .D(n958), .CLK(clk), .RSTB(n2373), .Q(reg29[15]) );
  DFFARX1 \regf_reg[28][14]  ( .D(n957), .CLK(clk), .RSTB(n2373), .Q(reg29[14]) );
  DFFARX1 \regf_reg[28][13]  ( .D(n956), .CLK(clk), .RSTB(n2373), .Q(reg29[13]) );
  DFFARX1 \regf_reg[28][12]  ( .D(n955), .CLK(clk), .RSTB(n2373), .Q(reg29[12]) );
  DFFARX1 \regf_reg[28][11]  ( .D(n954), .CLK(clk), .RSTB(n2372), .Q(reg29[11]) );
  DFFARX1 \regf_reg[28][10]  ( .D(n953), .CLK(clk), .RSTB(n2372), .Q(reg29[10]) );
  DFFARX1 \regf_reg[28][9]  ( .D(n952), .CLK(clk), .RSTB(n2372), .Q(reg29[9])
         );
  DFFARX1 \regf_reg[28][8]  ( .D(n951), .CLK(clk), .RSTB(n2372), .Q(reg29[8])
         );
  DFFARX1 \regf_reg[28][7]  ( .D(n950), .CLK(clk), .RSTB(n2372), .Q(reg29[7])
         );
  DFFARX1 \regf_reg[28][6]  ( .D(n949), .CLK(clk), .RSTB(n2372), .Q(reg29[6])
         );
  DFFARX1 \regf_reg[28][5]  ( .D(n948), .CLK(clk), .RSTB(n2372), .Q(reg29[5])
         );
  DFFARX1 \regf_reg[28][4]  ( .D(n947), .CLK(clk), .RSTB(n2372), .Q(reg29[4])
         );
  DFFARX1 \regf_reg[28][3]  ( .D(n946), .CLK(clk), .RSTB(n2372), .Q(reg29[3])
         );
  DFFARX1 \regf_reg[28][2]  ( .D(n945), .CLK(clk), .RSTB(n2372), .Q(reg29[2])
         );
  DFFARX1 \regf_reg[28][1]  ( .D(n944), .CLK(clk), .RSTB(n2372), .Q(reg29[1])
         );
  DFFARX1 \regf_reg[28][0]  ( .D(n943), .CLK(clk), .RSTB(n2372), .Q(reg29[0])
         );
  DFFARX1 \regf_reg[27][31]  ( .D(n942), .CLK(clk), .RSTB(n2371), .Q(reg28[31]) );
  DFFARX1 \regf_reg[27][30]  ( .D(n941), .CLK(clk), .RSTB(n2371), .Q(reg28[30]) );
  DFFARX1 \regf_reg[27][29]  ( .D(n940), .CLK(clk), .RSTB(n2371), .Q(reg28[29]) );
  DFFARX1 \regf_reg[27][28]  ( .D(n939), .CLK(clk), .RSTB(n2371), .Q(reg28[28]) );
  DFFARX1 \regf_reg[27][27]  ( .D(n938), .CLK(clk), .RSTB(n2371), .Q(reg28[27]) );
  DFFARX1 \regf_reg[27][26]  ( .D(n937), .CLK(clk), .RSTB(n2371), .Q(reg28[26]) );
  DFFARX1 \regf_reg[27][25]  ( .D(n936), .CLK(clk), .RSTB(n2371), .Q(reg28[25]) );
  DFFARX1 \regf_reg[27][24]  ( .D(n935), .CLK(clk), .RSTB(n2371), .Q(reg28[24]) );
  DFFARX1 \regf_reg[27][23]  ( .D(n934), .CLK(clk), .RSTB(n2371), .Q(reg28[23]) );
  DFFARX1 \regf_reg[27][22]  ( .D(n933), .CLK(clk), .RSTB(n2371), .Q(reg28[22]) );
  DFFARX1 \regf_reg[27][21]  ( .D(n932), .CLK(clk), .RSTB(n2371), .Q(reg28[21]) );
  DFFARX1 \regf_reg[27][20]  ( .D(n931), .CLK(clk), .RSTB(n2371), .Q(reg28[20]) );
  DFFARX1 \regf_reg[27][19]  ( .D(n930), .CLK(clk), .RSTB(n2370), .Q(reg28[19]) );
  DFFARX1 \regf_reg[27][18]  ( .D(n929), .CLK(clk), .RSTB(n2370), .Q(reg28[18]) );
  DFFARX1 \regf_reg[27][17]  ( .D(n928), .CLK(clk), .RSTB(n2370), .Q(reg28[17]) );
  DFFARX1 \regf_reg[27][16]  ( .D(n927), .CLK(clk), .RSTB(n2370), .Q(reg28[16]) );
  DFFARX1 \regf_reg[27][15]  ( .D(n926), .CLK(clk), .RSTB(n2370), .Q(reg28[15]) );
  DFFARX1 \regf_reg[27][14]  ( .D(n925), .CLK(clk), .RSTB(n2370), .Q(reg28[14]) );
  DFFARX1 \regf_reg[27][13]  ( .D(n924), .CLK(clk), .RSTB(n2370), .Q(reg28[13]) );
  DFFARX1 \regf_reg[27][12]  ( .D(n923), .CLK(clk), .RSTB(n2370), .Q(reg28[12]) );
  DFFARX1 \regf_reg[27][11]  ( .D(n922), .CLK(clk), .RSTB(n2370), .Q(reg28[11]) );
  DFFARX1 \regf_reg[27][10]  ( .D(n921), .CLK(clk), .RSTB(n2370), .Q(reg28[10]) );
  DFFARX1 \regf_reg[27][9]  ( .D(n920), .CLK(clk), .RSTB(n2370), .Q(reg28[9])
         );
  DFFARX1 \regf_reg[27][8]  ( .D(n919), .CLK(clk), .RSTB(n2370), .Q(reg28[8])
         );
  DFFARX1 \regf_reg[27][7]  ( .D(n918), .CLK(clk), .RSTB(n2369), .Q(reg28[7])
         );
  DFFARX1 \regf_reg[27][6]  ( .D(n917), .CLK(clk), .RSTB(n2369), .Q(reg28[6])
         );
  DFFARX1 \regf_reg[27][5]  ( .D(n916), .CLK(clk), .RSTB(n2369), .Q(reg28[5])
         );
  DFFARX1 \regf_reg[27][4]  ( .D(n915), .CLK(clk), .RSTB(n2369), .Q(reg28[4])
         );
  DFFARX1 \regf_reg[27][3]  ( .D(n914), .CLK(clk), .RSTB(n2369), .Q(reg28[3])
         );
  DFFARX1 \regf_reg[27][2]  ( .D(n913), .CLK(clk), .RSTB(n2369), .Q(reg28[2])
         );
  DFFARX1 \regf_reg[27][1]  ( .D(n912), .CLK(clk), .RSTB(n2369), .Q(reg28[1])
         );
  DFFARX1 \regf_reg[27][0]  ( .D(n911), .CLK(clk), .RSTB(n2369), .Q(reg28[0])
         );
  DFFARX1 \regf_reg[26][31]  ( .D(n910), .CLK(clk), .RSTB(n2369), .Q(reg27[31]) );
  DFFARX1 \regf_reg[26][30]  ( .D(n909), .CLK(clk), .RSTB(n2369), .Q(reg27[30]) );
  DFFARX1 \regf_reg[26][29]  ( .D(n908), .CLK(clk), .RSTB(n2369), .Q(reg27[29]) );
  DFFARX1 \regf_reg[26][28]  ( .D(n907), .CLK(clk), .RSTB(n2369), .Q(reg27[28]) );
  DFFARX1 \regf_reg[26][27]  ( .D(n906), .CLK(clk), .RSTB(n2368), .Q(reg27[27]) );
  DFFARX1 \regf_reg[26][26]  ( .D(n905), .CLK(clk), .RSTB(n2368), .Q(reg27[26]) );
  DFFARX1 \regf_reg[26][25]  ( .D(n904), .CLK(clk), .RSTB(n2368), .Q(reg27[25]) );
  DFFARX1 \regf_reg[26][24]  ( .D(n903), .CLK(clk), .RSTB(n2368), .Q(reg27[24]) );
  DFFARX1 \regf_reg[26][23]  ( .D(n902), .CLK(clk), .RSTB(n2368), .Q(reg27[23]) );
  DFFARX1 \regf_reg[26][22]  ( .D(n901), .CLK(clk), .RSTB(n2368), .Q(reg27[22]) );
  DFFARX1 \regf_reg[26][21]  ( .D(n900), .CLK(clk), .RSTB(n2368), .Q(reg27[21]) );
  DFFARX1 \regf_reg[26][20]  ( .D(n899), .CLK(clk), .RSTB(n2368), .Q(reg27[20]) );
  DFFARX1 \regf_reg[26][19]  ( .D(n898), .CLK(clk), .RSTB(n2368), .Q(reg27[19]) );
  DFFARX1 \regf_reg[26][18]  ( .D(n897), .CLK(clk), .RSTB(n2368), .Q(reg27[18]) );
  DFFARX1 \regf_reg[26][17]  ( .D(n896), .CLK(clk), .RSTB(n2368), .Q(reg27[17]) );
  DFFARX1 \regf_reg[26][16]  ( .D(n895), .CLK(clk), .RSTB(n2368), .Q(reg27[16]) );
  DFFARX1 \regf_reg[26][15]  ( .D(n894), .CLK(clk), .RSTB(n2367), .Q(reg27[15]) );
  DFFARX1 \regf_reg[26][14]  ( .D(n893), .CLK(clk), .RSTB(n2367), .Q(reg27[14]) );
  DFFARX1 \regf_reg[26][13]  ( .D(n892), .CLK(clk), .RSTB(n2367), .Q(reg27[13]) );
  DFFARX1 \regf_reg[26][12]  ( .D(n891), .CLK(clk), .RSTB(n2367), .Q(reg27[12]) );
  DFFARX1 \regf_reg[26][11]  ( .D(n890), .CLK(clk), .RSTB(n2367), .Q(reg27[11]) );
  DFFARX1 \regf_reg[26][10]  ( .D(n889), .CLK(clk), .RSTB(n2367), .Q(reg27[10]) );
  DFFARX1 \regf_reg[26][9]  ( .D(n888), .CLK(clk), .RSTB(n2367), .Q(reg27[9])
         );
  DFFARX1 \regf_reg[26][8]  ( .D(n887), .CLK(clk), .RSTB(n2367), .Q(reg27[8])
         );
  DFFARX1 \regf_reg[26][7]  ( .D(n886), .CLK(clk), .RSTB(n2367), .Q(reg27[7])
         );
  DFFARX1 \regf_reg[26][6]  ( .D(n885), .CLK(clk), .RSTB(n2367), .Q(reg27[6])
         );
  DFFARX1 \regf_reg[26][5]  ( .D(n884), .CLK(clk), .RSTB(n2367), .Q(reg27[5])
         );
  DFFARX1 \regf_reg[26][4]  ( .D(n883), .CLK(clk), .RSTB(n2367), .Q(reg27[4])
         );
  DFFARX1 \regf_reg[26][3]  ( .D(n882), .CLK(clk), .RSTB(n2366), .Q(reg27[3])
         );
  DFFARX1 \regf_reg[26][2]  ( .D(n881), .CLK(clk), .RSTB(n2366), .Q(reg27[2])
         );
  DFFARX1 \regf_reg[26][1]  ( .D(n880), .CLK(clk), .RSTB(n2366), .Q(reg27[1])
         );
  DFFARX1 \regf_reg[26][0]  ( .D(n879), .CLK(clk), .RSTB(n2366), .Q(reg27[0])
         );
  DFFARX1 \regf_reg[25][31]  ( .D(n878), .CLK(clk), .RSTB(n2366), .Q(reg26[31]) );
  DFFARX1 \regf_reg[25][30]  ( .D(n877), .CLK(clk), .RSTB(n2366), .Q(reg26[30]) );
  DFFARX1 \regf_reg[25][29]  ( .D(n876), .CLK(clk), .RSTB(n2366), .Q(reg26[29]) );
  DFFARX1 \regf_reg[25][28]  ( .D(n875), .CLK(clk), .RSTB(n2366), .Q(reg26[28]) );
  DFFARX1 \regf_reg[25][27]  ( .D(n874), .CLK(clk), .RSTB(n2366), .Q(reg26[27]) );
  DFFARX1 \regf_reg[25][26]  ( .D(n873), .CLK(clk), .RSTB(n2366), .Q(reg26[26]) );
  DFFARX1 \regf_reg[25][25]  ( .D(n872), .CLK(clk), .RSTB(n2366), .Q(reg26[25]) );
  DFFARX1 \regf_reg[25][24]  ( .D(n871), .CLK(clk), .RSTB(n2366), .Q(reg26[24]) );
  DFFARX1 \regf_reg[25][23]  ( .D(n870), .CLK(clk), .RSTB(n2365), .Q(reg26[23]) );
  DFFARX1 \regf_reg[25][22]  ( .D(n869), .CLK(clk), .RSTB(n2365), .Q(reg26[22]) );
  DFFARX1 \regf_reg[25][21]  ( .D(n868), .CLK(clk), .RSTB(n2365), .Q(reg26[21]) );
  DFFARX1 \regf_reg[25][20]  ( .D(n867), .CLK(clk), .RSTB(n2365), .Q(reg26[20]) );
  DFFARX1 \regf_reg[25][19]  ( .D(n866), .CLK(clk), .RSTB(n2365), .Q(reg26[19]) );
  DFFARX1 \regf_reg[25][18]  ( .D(n865), .CLK(clk), .RSTB(n2365), .Q(reg26[18]) );
  DFFARX1 \regf_reg[25][17]  ( .D(n864), .CLK(clk), .RSTB(n2365), .Q(reg26[17]) );
  DFFARX1 \regf_reg[25][16]  ( .D(n863), .CLK(clk), .RSTB(n2365), .Q(reg26[16]) );
  DFFARX1 \regf_reg[25][15]  ( .D(n862), .CLK(clk), .RSTB(n2365), .Q(reg26[15]) );
  DFFARX1 \regf_reg[25][14]  ( .D(n861), .CLK(clk), .RSTB(n2365), .Q(reg26[14]) );
  DFFARX1 \regf_reg[25][13]  ( .D(n860), .CLK(clk), .RSTB(n2365), .Q(reg26[13]) );
  DFFARX1 \regf_reg[25][12]  ( .D(n859), .CLK(clk), .RSTB(n2365), .Q(reg26[12]) );
  DFFARX1 \regf_reg[25][11]  ( .D(n858), .CLK(clk), .RSTB(n2364), .Q(reg26[11]) );
  DFFARX1 \regf_reg[25][10]  ( .D(n857), .CLK(clk), .RSTB(n2364), .Q(reg26[10]) );
  DFFARX1 \regf_reg[25][9]  ( .D(n856), .CLK(clk), .RSTB(n2364), .Q(reg26[9])
         );
  DFFARX1 \regf_reg[25][8]  ( .D(n855), .CLK(clk), .RSTB(n2364), .Q(reg26[8])
         );
  DFFARX1 \regf_reg[25][7]  ( .D(n854), .CLK(clk), .RSTB(n2364), .Q(reg26[7])
         );
  DFFARX1 \regf_reg[25][6]  ( .D(n853), .CLK(clk), .RSTB(n2364), .Q(reg26[6])
         );
  DFFARX1 \regf_reg[25][5]  ( .D(n852), .CLK(clk), .RSTB(n2364), .Q(reg26[5])
         );
  DFFARX1 \regf_reg[25][4]  ( .D(n851), .CLK(clk), .RSTB(n2364), .Q(reg26[4])
         );
  DFFARX1 \regf_reg[25][3]  ( .D(n850), .CLK(clk), .RSTB(n2364), .Q(reg26[3])
         );
  DFFARX1 \regf_reg[25][2]  ( .D(n849), .CLK(clk), .RSTB(n2364), .Q(reg26[2])
         );
  DFFARX1 \regf_reg[25][1]  ( .D(n848), .CLK(clk), .RSTB(n2364), .Q(reg26[1])
         );
  DFFARX1 \regf_reg[25][0]  ( .D(n847), .CLK(clk), .RSTB(n2364), .Q(reg26[0])
         );
  DFFARX1 \regf_reg[24][31]  ( .D(n846), .CLK(clk), .RSTB(n2363), .Q(reg25[31]) );
  DFFARX1 \regf_reg[24][30]  ( .D(n845), .CLK(clk), .RSTB(n2363), .Q(reg25[30]) );
  DFFARX1 \regf_reg[24][29]  ( .D(n844), .CLK(clk), .RSTB(n2363), .Q(reg25[29]) );
  DFFARX1 \regf_reg[24][28]  ( .D(n843), .CLK(clk), .RSTB(n2363), .Q(reg25[28]) );
  DFFARX1 \regf_reg[24][27]  ( .D(n842), .CLK(clk), .RSTB(n2363), .Q(reg25[27]) );
  DFFARX1 \regf_reg[24][26]  ( .D(n841), .CLK(clk), .RSTB(n2363), .Q(reg25[26]) );
  DFFARX1 \regf_reg[24][25]  ( .D(n840), .CLK(clk), .RSTB(n2363), .Q(reg25[25]) );
  DFFARX1 \regf_reg[24][24]  ( .D(n839), .CLK(clk), .RSTB(n2363), .Q(reg25[24]) );
  DFFARX1 \regf_reg[24][23]  ( .D(n838), .CLK(clk), .RSTB(n2363), .Q(reg25[23]) );
  DFFARX1 \regf_reg[24][22]  ( .D(n837), .CLK(clk), .RSTB(n2363), .Q(reg25[22]) );
  DFFARX1 \regf_reg[24][21]  ( .D(n836), .CLK(clk), .RSTB(n2363), .Q(reg25[21]) );
  DFFARX1 \regf_reg[24][20]  ( .D(n835), .CLK(clk), .RSTB(n2363), .Q(reg25[20]) );
  DFFARX1 \regf_reg[24][19]  ( .D(n834), .CLK(clk), .RSTB(n2362), .Q(reg25[19]) );
  DFFARX1 \regf_reg[24][18]  ( .D(n833), .CLK(clk), .RSTB(n2362), .Q(reg25[18]) );
  DFFARX1 \regf_reg[24][17]  ( .D(n832), .CLK(clk), .RSTB(n2362), .Q(reg25[17]) );
  DFFARX1 \regf_reg[24][16]  ( .D(n831), .CLK(clk), .RSTB(n2362), .Q(reg25[16]) );
  DFFARX1 \regf_reg[24][15]  ( .D(n830), .CLK(clk), .RSTB(n2362), .Q(reg25[15]) );
  DFFARX1 \regf_reg[24][14]  ( .D(n829), .CLK(clk), .RSTB(n2362), .Q(reg25[14]) );
  DFFARX1 \regf_reg[24][13]  ( .D(n828), .CLK(clk), .RSTB(n2362), .Q(reg25[13]) );
  DFFARX1 \regf_reg[24][12]  ( .D(n827), .CLK(clk), .RSTB(n2362), .Q(reg25[12]) );
  DFFARX1 \regf_reg[24][11]  ( .D(n826), .CLK(clk), .RSTB(n2362), .Q(reg25[11]) );
  DFFARX1 \regf_reg[24][10]  ( .D(n825), .CLK(clk), .RSTB(n2362), .Q(reg25[10]) );
  DFFARX1 \regf_reg[24][9]  ( .D(n824), .CLK(clk), .RSTB(n2362), .Q(reg25[9])
         );
  DFFARX1 \regf_reg[24][8]  ( .D(n823), .CLK(clk), .RSTB(n2362), .Q(reg25[8])
         );
  DFFARX1 \regf_reg[24][7]  ( .D(n822), .CLK(clk), .RSTB(n2361), .Q(reg25[7])
         );
  DFFARX1 \regf_reg[24][6]  ( .D(n821), .CLK(clk), .RSTB(n2361), .Q(reg25[6])
         );
  DFFARX1 \regf_reg[24][5]  ( .D(n820), .CLK(clk), .RSTB(n2361), .Q(reg25[5])
         );
  DFFARX1 \regf_reg[24][4]  ( .D(n819), .CLK(clk), .RSTB(n2361), .Q(reg25[4])
         );
  DFFARX1 \regf_reg[24][3]  ( .D(n818), .CLK(clk), .RSTB(n2361), .Q(reg25[3])
         );
  DFFARX1 \regf_reg[24][2]  ( .D(n817), .CLK(clk), .RSTB(n2361), .Q(reg25[2])
         );
  DFFARX1 \regf_reg[24][1]  ( .D(n816), .CLK(clk), .RSTB(n2361), .Q(reg25[1])
         );
  DFFARX1 \regf_reg[24][0]  ( .D(n815), .CLK(clk), .RSTB(n2361), .Q(reg25[0])
         );
  DFFARX1 \regf_reg[23][31]  ( .D(n814), .CLK(clk), .RSTB(n2361), .Q(reg24[31]) );
  DFFARX1 \regf_reg[23][30]  ( .D(n813), .CLK(clk), .RSTB(n2361), .Q(reg24[30]) );
  DFFARX1 \regf_reg[23][29]  ( .D(n812), .CLK(clk), .RSTB(n2361), .Q(reg24[29]) );
  DFFARX1 \regf_reg[23][28]  ( .D(n811), .CLK(clk), .RSTB(n2361), .Q(reg24[28]) );
  DFFARX1 \regf_reg[23][27]  ( .D(n810), .CLK(clk), .RSTB(n2360), .Q(reg24[27]) );
  DFFARX1 \regf_reg[23][26]  ( .D(n809), .CLK(clk), .RSTB(n2360), .Q(reg24[26]) );
  DFFARX1 \regf_reg[23][25]  ( .D(n808), .CLK(clk), .RSTB(n2360), .Q(reg24[25]) );
  DFFARX1 \regf_reg[23][24]  ( .D(n807), .CLK(clk), .RSTB(n2360), .Q(reg24[24]) );
  DFFARX1 \regf_reg[23][23]  ( .D(n806), .CLK(clk), .RSTB(n2360), .Q(reg24[23]) );
  DFFARX1 \regf_reg[23][22]  ( .D(n805), .CLK(clk), .RSTB(n2360), .Q(reg24[22]) );
  DFFARX1 \regf_reg[23][21]  ( .D(n804), .CLK(clk), .RSTB(n2360), .Q(reg24[21]) );
  DFFARX1 \regf_reg[23][20]  ( .D(n803), .CLK(clk), .RSTB(n2360), .Q(reg24[20]) );
  DFFARX1 \regf_reg[23][19]  ( .D(n802), .CLK(clk), .RSTB(n2360), .Q(reg24[19]) );
  DFFARX1 \regf_reg[23][18]  ( .D(n801), .CLK(clk), .RSTB(n2360), .Q(reg24[18]) );
  DFFARX1 \regf_reg[23][17]  ( .D(n800), .CLK(clk), .RSTB(n2360), .Q(reg24[17]) );
  DFFARX1 \regf_reg[23][16]  ( .D(n799), .CLK(clk), .RSTB(n2360), .Q(reg24[16]) );
  DFFARX1 \regf_reg[23][15]  ( .D(n798), .CLK(clk), .RSTB(n2359), .Q(reg24[15]) );
  DFFARX1 \regf_reg[23][14]  ( .D(n797), .CLK(clk), .RSTB(n2359), .Q(reg24[14]) );
  DFFARX1 \regf_reg[23][13]  ( .D(n796), .CLK(clk), .RSTB(n2359), .Q(reg24[13]) );
  DFFARX1 \regf_reg[23][12]  ( .D(n795), .CLK(clk), .RSTB(n2359), .Q(reg24[12]) );
  DFFARX1 \regf_reg[23][11]  ( .D(n794), .CLK(clk), .RSTB(n2359), .Q(reg24[11]) );
  DFFARX1 \regf_reg[23][10]  ( .D(n793), .CLK(clk), .RSTB(n2359), .Q(reg24[10]) );
  DFFARX1 \regf_reg[23][9]  ( .D(n792), .CLK(clk), .RSTB(n2359), .Q(reg24[9])
         );
  DFFARX1 \regf_reg[23][8]  ( .D(n791), .CLK(clk), .RSTB(n2359), .Q(reg24[8])
         );
  DFFARX1 \regf_reg[23][7]  ( .D(n790), .CLK(clk), .RSTB(n2359), .Q(reg24[7])
         );
  DFFARX1 \regf_reg[23][6]  ( .D(n789), .CLK(clk), .RSTB(n2359), .Q(reg24[6])
         );
  DFFARX1 \regf_reg[23][5]  ( .D(n788), .CLK(clk), .RSTB(n2359), .Q(reg24[5])
         );
  DFFARX1 \regf_reg[23][4]  ( .D(n787), .CLK(clk), .RSTB(n2359), .Q(reg24[4])
         );
  DFFARX1 \regf_reg[23][3]  ( .D(n786), .CLK(clk), .RSTB(n2358), .Q(reg24[3])
         );
  DFFARX1 \regf_reg[23][2]  ( .D(n785), .CLK(clk), .RSTB(n2358), .Q(reg24[2])
         );
  DFFARX1 \regf_reg[23][1]  ( .D(n784), .CLK(clk), .RSTB(n2358), .Q(reg24[1])
         );
  DFFARX1 \regf_reg[23][0]  ( .D(n783), .CLK(clk), .RSTB(n2358), .Q(reg24[0])
         );
  DFFARX1 \regf_reg[22][31]  ( .D(n782), .CLK(clk), .RSTB(n2358), .Q(reg23[31]) );
  DFFARX1 \regf_reg[22][30]  ( .D(n781), .CLK(clk), .RSTB(n2358), .Q(reg23[30]) );
  DFFARX1 \regf_reg[22][29]  ( .D(n780), .CLK(clk), .RSTB(n2358), .Q(reg23[29]) );
  DFFARX1 \regf_reg[22][28]  ( .D(n779), .CLK(clk), .RSTB(n2358), .Q(reg23[28]) );
  DFFARX1 \regf_reg[22][27]  ( .D(n778), .CLK(clk), .RSTB(n2358), .Q(reg23[27]) );
  DFFARX1 \regf_reg[22][26]  ( .D(n777), .CLK(clk), .RSTB(n2358), .Q(reg23[26]) );
  DFFARX1 \regf_reg[22][25]  ( .D(n776), .CLK(clk), .RSTB(n2358), .Q(reg23[25]) );
  DFFARX1 \regf_reg[22][24]  ( .D(n775), .CLK(clk), .RSTB(n2358), .Q(reg23[24]) );
  DFFARX1 \regf_reg[22][23]  ( .D(n774), .CLK(clk), .RSTB(n2357), .Q(reg23[23]) );
  DFFARX1 \regf_reg[22][22]  ( .D(n773), .CLK(clk), .RSTB(n2357), .Q(reg23[22]) );
  DFFARX1 \regf_reg[22][21]  ( .D(n772), .CLK(clk), .RSTB(n2357), .Q(reg23[21]) );
  DFFARX1 \regf_reg[22][20]  ( .D(n771), .CLK(clk), .RSTB(n2357), .Q(reg23[20]) );
  DFFARX1 \regf_reg[22][19]  ( .D(n770), .CLK(clk), .RSTB(n2357), .Q(reg23[19]) );
  DFFARX1 \regf_reg[22][18]  ( .D(n769), .CLK(clk), .RSTB(n2357), .Q(reg23[18]) );
  DFFARX1 \regf_reg[22][17]  ( .D(n768), .CLK(clk), .RSTB(n2357), .Q(reg23[17]) );
  DFFARX1 \regf_reg[22][16]  ( .D(n767), .CLK(clk), .RSTB(n2357), .Q(reg23[16]) );
  DFFARX1 \regf_reg[22][15]  ( .D(n766), .CLK(clk), .RSTB(n2357), .Q(reg23[15]) );
  DFFARX1 \regf_reg[22][14]  ( .D(n765), .CLK(clk), .RSTB(n2357), .Q(reg23[14]) );
  DFFARX1 \regf_reg[22][13]  ( .D(n764), .CLK(clk), .RSTB(n2357), .Q(reg23[13]) );
  DFFARX1 \regf_reg[22][12]  ( .D(n763), .CLK(clk), .RSTB(n2357), .Q(reg23[12]) );
  DFFARX1 \regf_reg[22][11]  ( .D(n762), .CLK(clk), .RSTB(n2356), .Q(reg23[11]) );
  DFFARX1 \regf_reg[22][10]  ( .D(n761), .CLK(clk), .RSTB(n2356), .Q(reg23[10]) );
  DFFARX1 \regf_reg[22][9]  ( .D(n760), .CLK(clk), .RSTB(n2356), .Q(reg23[9])
         );
  DFFARX1 \regf_reg[22][8]  ( .D(n759), .CLK(clk), .RSTB(n2356), .Q(reg23[8])
         );
  DFFARX1 \regf_reg[22][7]  ( .D(n758), .CLK(clk), .RSTB(n2356), .Q(reg23[7])
         );
  DFFARX1 \regf_reg[22][6]  ( .D(n757), .CLK(clk), .RSTB(n2356), .Q(reg23[6])
         );
  DFFARX1 \regf_reg[22][5]  ( .D(n756), .CLK(clk), .RSTB(n2356), .Q(reg23[5])
         );
  DFFARX1 \regf_reg[22][4]  ( .D(n755), .CLK(clk), .RSTB(n2356), .Q(reg23[4])
         );
  DFFARX1 \regf_reg[22][3]  ( .D(n754), .CLK(clk), .RSTB(n2356), .Q(reg23[3])
         );
  DFFARX1 \regf_reg[22][2]  ( .D(n753), .CLK(clk), .RSTB(n2356), .Q(reg23[2])
         );
  DFFARX1 \regf_reg[22][1]  ( .D(n752), .CLK(clk), .RSTB(n2356), .Q(reg23[1])
         );
  DFFARX1 \regf_reg[22][0]  ( .D(n751), .CLK(clk), .RSTB(n2356), .Q(reg23[0])
         );
  DFFARX1 \regf_reg[21][31]  ( .D(n750), .CLK(clk), .RSTB(n2355), .Q(reg22[31]) );
  DFFARX1 \regf_reg[21][30]  ( .D(n749), .CLK(clk), .RSTB(n2355), .Q(reg22[30]) );
  DFFARX1 \regf_reg[21][29]  ( .D(n748), .CLK(clk), .RSTB(n2355), .Q(reg22[29]) );
  DFFARX1 \regf_reg[21][28]  ( .D(n747), .CLK(clk), .RSTB(n2355), .Q(reg22[28]) );
  DFFARX1 \regf_reg[21][27]  ( .D(n746), .CLK(clk), .RSTB(n2355), .Q(reg22[27]) );
  DFFARX1 \regf_reg[21][26]  ( .D(n745), .CLK(clk), .RSTB(n2355), .Q(reg22[26]) );
  DFFARX1 \regf_reg[21][25]  ( .D(n744), .CLK(clk), .RSTB(n2355), .Q(reg22[25]) );
  DFFARX1 \regf_reg[21][24]  ( .D(n743), .CLK(clk), .RSTB(n2355), .Q(reg22[24]) );
  DFFARX1 \regf_reg[21][23]  ( .D(n742), .CLK(clk), .RSTB(n2355), .Q(reg22[23]) );
  DFFARX1 \regf_reg[21][22]  ( .D(n741), .CLK(clk), .RSTB(n2355), .Q(reg22[22]) );
  DFFARX1 \regf_reg[21][21]  ( .D(n740), .CLK(clk), .RSTB(n2355), .Q(reg22[21]) );
  DFFARX1 \regf_reg[21][20]  ( .D(n739), .CLK(clk), .RSTB(n2355), .Q(reg22[20]) );
  DFFARX1 \regf_reg[21][19]  ( .D(n738), .CLK(clk), .RSTB(n2354), .Q(reg22[19]) );
  DFFARX1 \regf_reg[21][18]  ( .D(n737), .CLK(clk), .RSTB(n2354), .Q(reg22[18]) );
  DFFARX1 \regf_reg[21][17]  ( .D(n736), .CLK(clk), .RSTB(n2354), .Q(reg22[17]) );
  DFFARX1 \regf_reg[21][16]  ( .D(n735), .CLK(clk), .RSTB(n2354), .Q(reg22[16]) );
  DFFARX1 \regf_reg[21][15]  ( .D(n734), .CLK(clk), .RSTB(n2354), .Q(reg22[15]) );
  DFFARX1 \regf_reg[21][14]  ( .D(n733), .CLK(clk), .RSTB(n2354), .Q(reg22[14]) );
  DFFARX1 \regf_reg[21][13]  ( .D(n732), .CLK(clk), .RSTB(n2354), .Q(reg22[13]) );
  DFFARX1 \regf_reg[21][12]  ( .D(n731), .CLK(clk), .RSTB(n2354), .Q(reg22[12]) );
  DFFARX1 \regf_reg[21][11]  ( .D(n730), .CLK(clk), .RSTB(n2354), .Q(reg22[11]) );
  DFFARX1 \regf_reg[21][10]  ( .D(n729), .CLK(clk), .RSTB(n2354), .Q(reg22[10]) );
  DFFARX1 \regf_reg[21][9]  ( .D(n728), .CLK(clk), .RSTB(n2354), .Q(reg22[9])
         );
  DFFARX1 \regf_reg[21][8]  ( .D(n727), .CLK(clk), .RSTB(n2354), .Q(reg22[8])
         );
  DFFARX1 \regf_reg[21][7]  ( .D(n726), .CLK(clk), .RSTB(n2353), .Q(reg22[7])
         );
  DFFARX1 \regf_reg[21][6]  ( .D(n725), .CLK(clk), .RSTB(n2353), .Q(reg22[6])
         );
  DFFARX1 \regf_reg[21][5]  ( .D(n724), .CLK(clk), .RSTB(n2353), .Q(reg22[5])
         );
  DFFARX1 \regf_reg[21][4]  ( .D(n723), .CLK(clk), .RSTB(n2353), .Q(reg22[4])
         );
  DFFARX1 \regf_reg[21][3]  ( .D(n722), .CLK(clk), .RSTB(n2353), .Q(reg22[3])
         );
  DFFARX1 \regf_reg[21][2]  ( .D(n721), .CLK(clk), .RSTB(n2353), .Q(reg22[2])
         );
  DFFARX1 \regf_reg[21][1]  ( .D(n720), .CLK(clk), .RSTB(n2353), .Q(reg22[1])
         );
  DFFARX1 \regf_reg[21][0]  ( .D(n719), .CLK(clk), .RSTB(n2353), .Q(reg22[0])
         );
  DFFARX1 \regf_reg[20][31]  ( .D(n718), .CLK(clk), .RSTB(n2353), .Q(reg21[31]) );
  DFFARX1 \regf_reg[20][30]  ( .D(n717), .CLK(clk), .RSTB(n2353), .Q(reg21[30]) );
  DFFARX1 \regf_reg[20][29]  ( .D(n716), .CLK(clk), .RSTB(n2353), .Q(reg21[29]) );
  DFFARX1 \regf_reg[20][28]  ( .D(n715), .CLK(clk), .RSTB(n2353), .Q(reg21[28]) );
  DFFARX1 \regf_reg[20][27]  ( .D(n714), .CLK(clk), .RSTB(n2352), .Q(reg21[27]) );
  DFFARX1 \regf_reg[20][26]  ( .D(n713), .CLK(clk), .RSTB(n2352), .Q(reg21[26]) );
  DFFARX1 \regf_reg[20][25]  ( .D(n712), .CLK(clk), .RSTB(n2352), .Q(reg21[25]) );
  DFFARX1 \regf_reg[20][24]  ( .D(n711), .CLK(clk), .RSTB(n2352), .Q(reg21[24]) );
  DFFARX1 \regf_reg[20][23]  ( .D(n710), .CLK(clk), .RSTB(n2352), .Q(reg21[23]) );
  DFFARX1 \regf_reg[20][22]  ( .D(n709), .CLK(clk), .RSTB(n2352), .Q(reg21[22]) );
  DFFARX1 \regf_reg[20][21]  ( .D(n708), .CLK(clk), .RSTB(n2352), .Q(reg21[21]) );
  DFFARX1 \regf_reg[20][20]  ( .D(n707), .CLK(clk), .RSTB(n2352), .Q(reg21[20]) );
  DFFARX1 \regf_reg[20][19]  ( .D(n706), .CLK(clk), .RSTB(n2352), .Q(reg21[19]) );
  DFFARX1 \regf_reg[20][18]  ( .D(n705), .CLK(clk), .RSTB(n2352), .Q(reg21[18]) );
  DFFARX1 \regf_reg[20][17]  ( .D(n704), .CLK(clk), .RSTB(n2352), .Q(reg21[17]) );
  DFFARX1 \regf_reg[20][16]  ( .D(n703), .CLK(clk), .RSTB(n2352), .Q(reg21[16]) );
  DFFARX1 \regf_reg[20][15]  ( .D(n702), .CLK(clk), .RSTB(n2351), .Q(reg21[15]) );
  DFFARX1 \regf_reg[20][14]  ( .D(n701), .CLK(clk), .RSTB(n2351), .Q(reg21[14]) );
  DFFARX1 \regf_reg[20][13]  ( .D(n700), .CLK(clk), .RSTB(n2351), .Q(reg21[13]) );
  DFFARX1 \regf_reg[20][12]  ( .D(n699), .CLK(clk), .RSTB(n2351), .Q(reg21[12]) );
  DFFARX1 \regf_reg[20][11]  ( .D(n698), .CLK(clk), .RSTB(n2351), .Q(reg21[11]) );
  DFFARX1 \regf_reg[20][10]  ( .D(n697), .CLK(clk), .RSTB(n2351), .Q(reg21[10]) );
  DFFARX1 \regf_reg[20][9]  ( .D(n696), .CLK(clk), .RSTB(n2351), .Q(reg21[9])
         );
  DFFARX1 \regf_reg[20][8]  ( .D(n695), .CLK(clk), .RSTB(n2351), .Q(reg21[8])
         );
  DFFARX1 \regf_reg[20][7]  ( .D(n694), .CLK(clk), .RSTB(n2351), .Q(reg21[7])
         );
  DFFARX1 \regf_reg[20][6]  ( .D(n693), .CLK(clk), .RSTB(n2351), .Q(reg21[6])
         );
  DFFARX1 \regf_reg[20][5]  ( .D(n692), .CLK(clk), .RSTB(n2351), .Q(reg21[5])
         );
  DFFARX1 \regf_reg[20][4]  ( .D(n691), .CLK(clk), .RSTB(n2351), .Q(reg21[4])
         );
  DFFARX1 \regf_reg[20][3]  ( .D(n690), .CLK(clk), .RSTB(n2350), .Q(reg21[3])
         );
  DFFARX1 \regf_reg[20][2]  ( .D(n689), .CLK(clk), .RSTB(n2350), .Q(reg21[2])
         );
  DFFARX1 \regf_reg[20][1]  ( .D(n688), .CLK(clk), .RSTB(n2350), .Q(reg21[1])
         );
  DFFARX1 \regf_reg[20][0]  ( .D(n687), .CLK(clk), .RSTB(n2350), .Q(reg21[0])
         );
  DFFARX1 \regf_reg[19][31]  ( .D(n686), .CLK(clk), .RSTB(n2350), .Q(reg20[31]) );
  DFFARX1 \regf_reg[19][30]  ( .D(n685), .CLK(clk), .RSTB(n2350), .Q(reg20[30]) );
  DFFARX1 \regf_reg[19][29]  ( .D(n684), .CLK(clk), .RSTB(n2350), .Q(reg20[29]) );
  DFFARX1 \regf_reg[19][28]  ( .D(n683), .CLK(clk), .RSTB(n2350), .Q(reg20[28]) );
  DFFARX1 \regf_reg[19][27]  ( .D(n682), .CLK(clk), .RSTB(n2350), .Q(reg20[27]) );
  DFFARX1 \regf_reg[19][26]  ( .D(n681), .CLK(clk), .RSTB(n2350), .Q(reg20[26]) );
  DFFARX1 \regf_reg[19][25]  ( .D(n680), .CLK(clk), .RSTB(n2350), .Q(reg20[25]) );
  DFFARX1 \regf_reg[19][24]  ( .D(n679), .CLK(clk), .RSTB(n2350), .Q(reg20[24]) );
  DFFARX1 \regf_reg[19][23]  ( .D(n678), .CLK(clk), .RSTB(n2349), .Q(reg20[23]) );
  DFFARX1 \regf_reg[19][22]  ( .D(n677), .CLK(clk), .RSTB(n2349), .Q(reg20[22]) );
  DFFARX1 \regf_reg[19][21]  ( .D(n676), .CLK(clk), .RSTB(n2349), .Q(reg20[21]) );
  DFFARX1 \regf_reg[19][20]  ( .D(n675), .CLK(clk), .RSTB(n2349), .Q(reg20[20]) );
  DFFARX1 \regf_reg[19][19]  ( .D(n674), .CLK(clk), .RSTB(n2349), .Q(reg20[19]) );
  DFFARX1 \regf_reg[19][18]  ( .D(n673), .CLK(clk), .RSTB(n2349), .Q(reg20[18]) );
  DFFARX1 \regf_reg[19][17]  ( .D(n672), .CLK(clk), .RSTB(n2349), .Q(reg20[17]) );
  DFFARX1 \regf_reg[19][16]  ( .D(n671), .CLK(clk), .RSTB(n2349), .Q(reg20[16]) );
  DFFARX1 \regf_reg[19][15]  ( .D(n670), .CLK(clk), .RSTB(n2349), .Q(reg20[15]) );
  DFFARX1 \regf_reg[19][14]  ( .D(n669), .CLK(clk), .RSTB(n2349), .Q(reg20[14]) );
  DFFARX1 \regf_reg[19][13]  ( .D(n668), .CLK(clk), .RSTB(n2349), .Q(reg20[13]) );
  DFFARX1 \regf_reg[19][12]  ( .D(n667), .CLK(clk), .RSTB(n2349), .Q(reg20[12]) );
  DFFARX1 \regf_reg[19][11]  ( .D(n666), .CLK(clk), .RSTB(n2348), .Q(reg20[11]) );
  DFFARX1 \regf_reg[19][10]  ( .D(n665), .CLK(clk), .RSTB(n2348), .Q(reg20[10]) );
  DFFARX1 \regf_reg[19][9]  ( .D(n664), .CLK(clk), .RSTB(n2348), .Q(reg20[9])
         );
  DFFARX1 \regf_reg[19][8]  ( .D(n663), .CLK(clk), .RSTB(n2348), .Q(reg20[8])
         );
  DFFARX1 \regf_reg[19][7]  ( .D(n662), .CLK(clk), .RSTB(n2348), .Q(reg20[7])
         );
  DFFARX1 \regf_reg[19][6]  ( .D(n661), .CLK(clk), .RSTB(n2348), .Q(reg20[6])
         );
  DFFARX1 \regf_reg[19][5]  ( .D(n660), .CLK(clk), .RSTB(n2348), .Q(reg20[5])
         );
  DFFARX1 \regf_reg[19][4]  ( .D(n659), .CLK(clk), .RSTB(n2348), .Q(reg20[4])
         );
  DFFARX1 \regf_reg[19][3]  ( .D(n658), .CLK(clk), .RSTB(n2348), .Q(reg20[3])
         );
  DFFARX1 \regf_reg[19][2]  ( .D(n657), .CLK(clk), .RSTB(n2348), .Q(reg20[2])
         );
  DFFARX1 \regf_reg[19][1]  ( .D(n656), .CLK(clk), .RSTB(n2348), .Q(reg20[1])
         );
  DFFARX1 \regf_reg[19][0]  ( .D(n655), .CLK(clk), .RSTB(n2348), .Q(reg20[0])
         );
  DFFARX1 \regf_reg[18][31]  ( .D(n654), .CLK(clk), .RSTB(n2347), .Q(reg19[31]) );
  DFFARX1 \regf_reg[18][30]  ( .D(n653), .CLK(clk), .RSTB(n2347), .Q(reg19[30]) );
  DFFARX1 \regf_reg[18][29]  ( .D(n652), .CLK(clk), .RSTB(n2347), .Q(reg19[29]) );
  DFFARX1 \regf_reg[18][28]  ( .D(n651), .CLK(clk), .RSTB(n2347), .Q(reg19[28]) );
  DFFARX1 \regf_reg[18][27]  ( .D(n650), .CLK(clk), .RSTB(n2347), .Q(reg19[27]) );
  DFFARX1 \regf_reg[18][26]  ( .D(n649), .CLK(clk), .RSTB(n2347), .Q(reg19[26]) );
  DFFARX1 \regf_reg[18][25]  ( .D(n648), .CLK(clk), .RSTB(n2347), .Q(reg19[25]) );
  DFFARX1 \regf_reg[18][24]  ( .D(n647), .CLK(clk), .RSTB(n2347), .Q(reg19[24]) );
  DFFARX1 \regf_reg[18][23]  ( .D(n646), .CLK(clk), .RSTB(n2347), .Q(reg19[23]) );
  DFFARX1 \regf_reg[18][22]  ( .D(n645), .CLK(clk), .RSTB(n2347), .Q(reg19[22]) );
  DFFARX1 \regf_reg[18][21]  ( .D(n644), .CLK(clk), .RSTB(n2347), .Q(reg19[21]) );
  DFFARX1 \regf_reg[18][20]  ( .D(n643), .CLK(clk), .RSTB(n2347), .Q(reg19[20]) );
  DFFARX1 \regf_reg[18][19]  ( .D(n642), .CLK(clk), .RSTB(n2346), .Q(reg19[19]) );
  DFFARX1 \regf_reg[18][18]  ( .D(n641), .CLK(clk), .RSTB(n2346), .Q(reg19[18]) );
  DFFARX1 \regf_reg[18][17]  ( .D(n640), .CLK(clk), .RSTB(n2346), .Q(reg19[17]) );
  DFFARX1 \regf_reg[18][16]  ( .D(n639), .CLK(clk), .RSTB(n2346), .Q(reg19[16]) );
  DFFARX1 \regf_reg[18][15]  ( .D(n638), .CLK(clk), .RSTB(n2346), .Q(reg19[15]) );
  DFFARX1 \regf_reg[18][14]  ( .D(n637), .CLK(clk), .RSTB(n2346), .Q(reg19[14]) );
  DFFARX1 \regf_reg[18][13]  ( .D(n636), .CLK(clk), .RSTB(n2346), .Q(reg19[13]) );
  DFFARX1 \regf_reg[18][12]  ( .D(n635), .CLK(clk), .RSTB(n2346), .Q(reg19[12]) );
  DFFARX1 \regf_reg[18][11]  ( .D(n634), .CLK(clk), .RSTB(n2346), .Q(reg19[11]) );
  DFFARX1 \regf_reg[18][10]  ( .D(n633), .CLK(clk), .RSTB(n2346), .Q(reg19[10]) );
  DFFARX1 \regf_reg[18][9]  ( .D(n632), .CLK(clk), .RSTB(n2346), .Q(reg19[9])
         );
  DFFARX1 \regf_reg[18][8]  ( .D(n631), .CLK(clk), .RSTB(n2346), .Q(reg19[8])
         );
  DFFARX1 \regf_reg[18][7]  ( .D(n630), .CLK(clk), .RSTB(n2345), .Q(reg19[7])
         );
  DFFARX1 \regf_reg[18][6]  ( .D(n629), .CLK(clk), .RSTB(n2345), .Q(reg19[6])
         );
  DFFARX1 \regf_reg[18][5]  ( .D(n628), .CLK(clk), .RSTB(n2345), .Q(reg19[5])
         );
  DFFARX1 \regf_reg[18][4]  ( .D(n627), .CLK(clk), .RSTB(n2345), .Q(reg19[4])
         );
  DFFARX1 \regf_reg[18][3]  ( .D(n626), .CLK(clk), .RSTB(n2345), .Q(reg19[3])
         );
  DFFARX1 \regf_reg[18][2]  ( .D(n625), .CLK(clk), .RSTB(n2345), .Q(reg19[2])
         );
  DFFARX1 \regf_reg[18][1]  ( .D(n624), .CLK(clk), .RSTB(n2345), .Q(reg19[1])
         );
  DFFARX1 \regf_reg[18][0]  ( .D(n623), .CLK(clk), .RSTB(n2345), .Q(reg19[0])
         );
  DFFARX1 \regf_reg[17][31]  ( .D(n622), .CLK(clk), .RSTB(n2345), .Q(reg18[31]) );
  DFFARX1 \regf_reg[17][30]  ( .D(n621), .CLK(clk), .RSTB(n2345), .Q(reg18[30]) );
  DFFARX1 \regf_reg[17][29]  ( .D(n620), .CLK(clk), .RSTB(n2345), .Q(reg18[29]) );
  DFFARX1 \regf_reg[17][28]  ( .D(n619), .CLK(clk), .RSTB(n2345), .Q(reg18[28]) );
  DFFARX1 \regf_reg[17][27]  ( .D(n618), .CLK(clk), .RSTB(n2344), .Q(reg18[27]) );
  DFFARX1 \regf_reg[17][26]  ( .D(n617), .CLK(clk), .RSTB(n2344), .Q(reg18[26]) );
  DFFARX1 \regf_reg[17][25]  ( .D(n616), .CLK(clk), .RSTB(n2344), .Q(reg18[25]) );
  DFFARX1 \regf_reg[17][24]  ( .D(n615), .CLK(clk), .RSTB(n2344), .Q(reg18[24]) );
  DFFARX1 \regf_reg[17][23]  ( .D(n614), .CLK(clk), .RSTB(n2344), .Q(reg18[23]) );
  DFFARX1 \regf_reg[17][22]  ( .D(n613), .CLK(clk), .RSTB(n2344), .Q(reg18[22]) );
  DFFARX1 \regf_reg[17][21]  ( .D(n612), .CLK(clk), .RSTB(n2344), .Q(reg18[21]) );
  DFFARX1 \regf_reg[17][20]  ( .D(n611), .CLK(clk), .RSTB(n2344), .Q(reg18[20]) );
  DFFARX1 \regf_reg[17][19]  ( .D(n610), .CLK(clk), .RSTB(n2344), .Q(reg18[19]) );
  DFFARX1 \regf_reg[17][18]  ( .D(n609), .CLK(clk), .RSTB(n2344), .Q(reg18[18]) );
  DFFARX1 \regf_reg[17][17]  ( .D(n608), .CLK(clk), .RSTB(n2344), .Q(reg18[17]) );
  DFFARX1 \regf_reg[17][16]  ( .D(n607), .CLK(clk), .RSTB(n2344), .Q(reg18[16]) );
  DFFARX1 \regf_reg[17][15]  ( .D(n606), .CLK(clk), .RSTB(n2343), .Q(reg18[15]) );
  DFFARX1 \regf_reg[17][14]  ( .D(n605), .CLK(clk), .RSTB(n2343), .Q(reg18[14]) );
  DFFARX1 \regf_reg[17][13]  ( .D(n604), .CLK(clk), .RSTB(n2343), .Q(reg18[13]) );
  DFFARX1 \regf_reg[17][12]  ( .D(n603), .CLK(clk), .RSTB(n2343), .Q(reg18[12]) );
  DFFARX1 \regf_reg[17][11]  ( .D(n602), .CLK(clk), .RSTB(n2343), .Q(reg18[11]) );
  DFFARX1 \regf_reg[17][10]  ( .D(n601), .CLK(clk), .RSTB(n2343), .Q(reg18[10]) );
  DFFARX1 \regf_reg[17][9]  ( .D(n600), .CLK(clk), .RSTB(n2343), .Q(reg18[9])
         );
  DFFARX1 \regf_reg[17][8]  ( .D(n599), .CLK(clk), .RSTB(n2343), .Q(reg18[8])
         );
  DFFARX1 \regf_reg[17][7]  ( .D(n598), .CLK(clk), .RSTB(n2343), .Q(reg18[7])
         );
  DFFARX1 \regf_reg[17][6]  ( .D(n597), .CLK(clk), .RSTB(n2343), .Q(reg18[6])
         );
  DFFARX1 \regf_reg[17][5]  ( .D(n596), .CLK(clk), .RSTB(n2343), .Q(reg18[5])
         );
  DFFARX1 \regf_reg[17][4]  ( .D(n595), .CLK(clk), .RSTB(n2343), .Q(reg18[4])
         );
  DFFARX1 \regf_reg[17][3]  ( .D(n594), .CLK(clk), .RSTB(n2342), .Q(reg18[3])
         );
  DFFARX1 \regf_reg[17][2]  ( .D(n593), .CLK(clk), .RSTB(n2342), .Q(reg18[2])
         );
  DFFARX1 \regf_reg[17][1]  ( .D(n592), .CLK(clk), .RSTB(n2342), .Q(reg18[1])
         );
  DFFARX1 \regf_reg[17][0]  ( .D(n591), .CLK(clk), .RSTB(n2342), .Q(reg18[0])
         );
  DFFARX1 \regf_reg[16][31]  ( .D(n590), .CLK(clk), .RSTB(n2342), .Q(reg17[31]) );
  DFFARX1 \regf_reg[16][30]  ( .D(n589), .CLK(clk), .RSTB(n2342), .Q(reg17[30]) );
  DFFARX1 \regf_reg[16][29]  ( .D(n588), .CLK(clk), .RSTB(n2342), .Q(reg17[29]) );
  DFFARX1 \regf_reg[16][28]  ( .D(n587), .CLK(clk), .RSTB(n2342), .Q(reg17[28]) );
  DFFARX1 \regf_reg[16][27]  ( .D(n586), .CLK(clk), .RSTB(n2342), .Q(reg17[27]) );
  DFFARX1 \regf_reg[16][26]  ( .D(n585), .CLK(clk), .RSTB(n2342), .Q(reg17[26]) );
  DFFARX1 \regf_reg[16][25]  ( .D(n584), .CLK(clk), .RSTB(n2342), .Q(reg17[25]) );
  DFFARX1 \regf_reg[16][24]  ( .D(n583), .CLK(clk), .RSTB(n2342), .Q(reg17[24]) );
  DFFARX1 \regf_reg[16][23]  ( .D(n582), .CLK(clk), .RSTB(n2341), .Q(reg17[23]) );
  DFFARX1 \regf_reg[16][22]  ( .D(n581), .CLK(clk), .RSTB(n2341), .Q(reg17[22]) );
  DFFARX1 \regf_reg[16][21]  ( .D(n580), .CLK(clk), .RSTB(n2341), .Q(reg17[21]) );
  DFFARX1 \regf_reg[16][20]  ( .D(n579), .CLK(clk), .RSTB(n2341), .Q(reg17[20]) );
  DFFARX1 \regf_reg[16][19]  ( .D(n578), .CLK(clk), .RSTB(n2341), .Q(reg17[19]) );
  DFFARX1 \regf_reg[16][18]  ( .D(n577), .CLK(clk), .RSTB(n2341), .Q(reg17[18]) );
  DFFARX1 \regf_reg[16][17]  ( .D(n576), .CLK(clk), .RSTB(n2341), .Q(reg17[17]) );
  DFFARX1 \regf_reg[16][16]  ( .D(n575), .CLK(clk), .RSTB(n2341), .Q(reg17[16]) );
  DFFARX1 \regf_reg[16][15]  ( .D(n574), .CLK(clk), .RSTB(n2341), .Q(reg17[15]) );
  DFFARX1 \regf_reg[16][14]  ( .D(n573), .CLK(clk), .RSTB(n2341), .Q(reg17[14]) );
  DFFARX1 \regf_reg[16][13]  ( .D(n572), .CLK(clk), .RSTB(n2341), .Q(reg17[13]) );
  DFFARX1 \regf_reg[16][12]  ( .D(n571), .CLK(clk), .RSTB(n2341), .Q(reg17[12]) );
  DFFARX1 \regf_reg[16][11]  ( .D(n570), .CLK(clk), .RSTB(n2340), .Q(reg17[11]) );
  DFFARX1 \regf_reg[16][10]  ( .D(n569), .CLK(clk), .RSTB(n2340), .Q(reg17[10]) );
  DFFARX1 \regf_reg[16][9]  ( .D(n568), .CLK(clk), .RSTB(n2340), .Q(reg17[9])
         );
  DFFARX1 \regf_reg[16][8]  ( .D(n567), .CLK(clk), .RSTB(n2340), .Q(reg17[8])
         );
  DFFARX1 \regf_reg[16][7]  ( .D(n566), .CLK(clk), .RSTB(n2340), .Q(reg17[7])
         );
  DFFARX1 \regf_reg[16][6]  ( .D(n565), .CLK(clk), .RSTB(n2340), .Q(reg17[6])
         );
  DFFARX1 \regf_reg[16][5]  ( .D(n564), .CLK(clk), .RSTB(n2340), .Q(reg17[5])
         );
  DFFARX1 \regf_reg[16][4]  ( .D(n563), .CLK(clk), .RSTB(n2340), .Q(reg17[4])
         );
  DFFARX1 \regf_reg[16][3]  ( .D(n562), .CLK(clk), .RSTB(n2340), .Q(reg17[3])
         );
  DFFARX1 \regf_reg[16][2]  ( .D(n561), .CLK(clk), .RSTB(n2340), .Q(reg17[2])
         );
  DFFARX1 \regf_reg[16][1]  ( .D(n560), .CLK(clk), .RSTB(n2340), .Q(reg17[1])
         );
  DFFARX1 \regf_reg[16][0]  ( .D(n559), .CLK(clk), .RSTB(n2340), .Q(reg17[0])
         );
  DFFARX1 \regf_reg[15][31]  ( .D(n558), .CLK(clk), .RSTB(n2339), .Q(reg16[31]) );
  DFFARX1 \regf_reg[15][30]  ( .D(n557), .CLK(clk), .RSTB(n2339), .Q(reg16[30]) );
  DFFARX1 \regf_reg[15][29]  ( .D(n556), .CLK(clk), .RSTB(n2339), .Q(reg16[29]) );
  DFFARX1 \regf_reg[15][28]  ( .D(n555), .CLK(clk), .RSTB(n2339), .Q(reg16[28]) );
  DFFARX1 \regf_reg[15][27]  ( .D(n554), .CLK(clk), .RSTB(n2339), .Q(reg16[27]) );
  DFFARX1 \regf_reg[15][26]  ( .D(n553), .CLK(clk), .RSTB(n2339), .Q(reg16[26]) );
  DFFARX1 \regf_reg[15][25]  ( .D(n552), .CLK(clk), .RSTB(n2339), .Q(reg16[25]) );
  DFFARX1 \regf_reg[15][24]  ( .D(n551), .CLK(clk), .RSTB(n2339), .Q(reg16[24]) );
  DFFARX1 \regf_reg[15][23]  ( .D(n550), .CLK(clk), .RSTB(n2339), .Q(reg16[23]) );
  DFFARX1 \regf_reg[15][22]  ( .D(n549), .CLK(clk), .RSTB(n2339), .Q(reg16[22]) );
  DFFARX1 \regf_reg[15][21]  ( .D(n548), .CLK(clk), .RSTB(n2339), .Q(reg16[21]) );
  DFFARX1 \regf_reg[15][20]  ( .D(n547), .CLK(clk), .RSTB(n2339), .Q(reg16[20]) );
  DFFARX1 \regf_reg[15][19]  ( .D(n546), .CLK(clk), .RSTB(n2338), .Q(reg16[19]) );
  DFFARX1 \regf_reg[15][18]  ( .D(n545), .CLK(clk), .RSTB(n2338), .Q(reg16[18]) );
  DFFARX1 \regf_reg[15][17]  ( .D(n544), .CLK(clk), .RSTB(n2338), .Q(reg16[17]) );
  DFFARX1 \regf_reg[15][16]  ( .D(n543), .CLK(clk), .RSTB(n2338), .Q(reg16[16]) );
  DFFARX1 \regf_reg[15][15]  ( .D(n542), .CLK(clk), .RSTB(n2338), .Q(reg16[15]) );
  DFFARX1 \regf_reg[15][14]  ( .D(n541), .CLK(clk), .RSTB(n2338), .Q(reg16[14]) );
  DFFARX1 \regf_reg[15][13]  ( .D(n540), .CLK(clk), .RSTB(n2338), .Q(reg16[13]) );
  DFFARX1 \regf_reg[15][12]  ( .D(n539), .CLK(clk), .RSTB(n2338), .Q(reg16[12]) );
  DFFARX1 \regf_reg[15][11]  ( .D(n538), .CLK(clk), .RSTB(n2338), .Q(reg16[11]) );
  DFFARX1 \regf_reg[15][10]  ( .D(n537), .CLK(clk), .RSTB(n2338), .Q(reg16[10]) );
  DFFARX1 \regf_reg[15][9]  ( .D(n536), .CLK(clk), .RSTB(n2338), .Q(reg16[9])
         );
  DFFARX1 \regf_reg[15][8]  ( .D(n535), .CLK(clk), .RSTB(n2338), .Q(reg16[8])
         );
  DFFARX1 \regf_reg[15][7]  ( .D(n534), .CLK(clk), .RSTB(n2337), .Q(reg16[7])
         );
  DFFARX1 \regf_reg[15][6]  ( .D(n533), .CLK(clk), .RSTB(n2337), .Q(reg16[6])
         );
  DFFARX1 \regf_reg[15][5]  ( .D(n532), .CLK(clk), .RSTB(n2337), .Q(reg16[5])
         );
  DFFARX1 \regf_reg[15][4]  ( .D(n531), .CLK(clk), .RSTB(n2337), .Q(reg16[4])
         );
  DFFARX1 \regf_reg[15][3]  ( .D(n530), .CLK(clk), .RSTB(n2337), .Q(reg16[3])
         );
  DFFARX1 \regf_reg[15][2]  ( .D(n529), .CLK(clk), .RSTB(n2337), .Q(reg16[2])
         );
  DFFARX1 \regf_reg[15][1]  ( .D(n528), .CLK(clk), .RSTB(n2337), .Q(reg16[1])
         );
  DFFARX1 \regf_reg[15][0]  ( .D(n527), .CLK(clk), .RSTB(n2337), .Q(reg16[0])
         );
  DFFARX1 \regf_reg[14][31]  ( .D(n526), .CLK(clk), .RSTB(n2337), .Q(reg15[31]) );
  DFFARX1 \regf_reg[14][30]  ( .D(n525), .CLK(clk), .RSTB(n2337), .Q(reg15[30]) );
  DFFARX1 \regf_reg[14][29]  ( .D(n524), .CLK(clk), .RSTB(n2337), .Q(reg15[29]) );
  DFFARX1 \regf_reg[14][28]  ( .D(n523), .CLK(clk), .RSTB(n2337), .Q(reg15[28]) );
  DFFARX1 \regf_reg[14][27]  ( .D(n522), .CLK(clk), .RSTB(n2336), .Q(reg15[27]) );
  DFFARX1 \regf_reg[14][26]  ( .D(n521), .CLK(clk), .RSTB(n2336), .Q(reg15[26]) );
  DFFARX1 \regf_reg[14][25]  ( .D(n520), .CLK(clk), .RSTB(n2336), .Q(reg15[25]) );
  DFFARX1 \regf_reg[14][24]  ( .D(n519), .CLK(clk), .RSTB(n2336), .Q(reg15[24]) );
  DFFARX1 \regf_reg[14][23]  ( .D(n518), .CLK(clk), .RSTB(n2336), .Q(reg15[23]) );
  DFFARX1 \regf_reg[14][22]  ( .D(n517), .CLK(clk), .RSTB(n2336), .Q(reg15[22]) );
  DFFARX1 \regf_reg[14][21]  ( .D(n516), .CLK(clk), .RSTB(n2336), .Q(reg15[21]) );
  DFFARX1 \regf_reg[14][20]  ( .D(n515), .CLK(clk), .RSTB(n2336), .Q(reg15[20]) );
  DFFARX1 \regf_reg[14][19]  ( .D(n514), .CLK(clk), .RSTB(n2336), .Q(reg15[19]) );
  DFFARX1 \regf_reg[14][18]  ( .D(n513), .CLK(clk), .RSTB(n2336), .Q(reg15[18]) );
  DFFARX1 \regf_reg[14][17]  ( .D(n512), .CLK(clk), .RSTB(n2336), .Q(reg15[17]) );
  DFFARX1 \regf_reg[14][16]  ( .D(n511), .CLK(clk), .RSTB(n2336), .Q(reg15[16]) );
  DFFARX1 \regf_reg[14][15]  ( .D(n510), .CLK(clk), .RSTB(n2335), .Q(reg15[15]) );
  DFFARX1 \regf_reg[14][14]  ( .D(n509), .CLK(clk), .RSTB(n2335), .Q(reg15[14]) );
  DFFARX1 \regf_reg[14][13]  ( .D(n508), .CLK(clk), .RSTB(n2335), .Q(reg15[13]) );
  DFFARX1 \regf_reg[14][12]  ( .D(n507), .CLK(clk), .RSTB(n2335), .Q(reg15[12]) );
  DFFARX1 \regf_reg[14][11]  ( .D(n506), .CLK(clk), .RSTB(n2335), .Q(reg15[11]) );
  DFFARX1 \regf_reg[14][10]  ( .D(n505), .CLK(clk), .RSTB(n2335), .Q(reg15[10]) );
  DFFARX1 \regf_reg[14][9]  ( .D(n504), .CLK(clk), .RSTB(n2335), .Q(reg15[9])
         );
  DFFARX1 \regf_reg[14][8]  ( .D(n503), .CLK(clk), .RSTB(n2335), .Q(reg15[8])
         );
  DFFARX1 \regf_reg[14][7]  ( .D(n502), .CLK(clk), .RSTB(n2335), .Q(reg15[7])
         );
  DFFARX1 \regf_reg[14][6]  ( .D(n501), .CLK(clk), .RSTB(n2335), .Q(reg15[6])
         );
  DFFARX1 \regf_reg[14][5]  ( .D(n500), .CLK(clk), .RSTB(n2335), .Q(reg15[5])
         );
  DFFARX1 \regf_reg[14][4]  ( .D(n499), .CLK(clk), .RSTB(n2335), .Q(reg15[4])
         );
  DFFARX1 \regf_reg[14][3]  ( .D(n498), .CLK(clk), .RSTB(n2334), .Q(reg15[3])
         );
  DFFARX1 \regf_reg[14][2]  ( .D(n497), .CLK(clk), .RSTB(n2334), .Q(reg15[2])
         );
  DFFARX1 \regf_reg[14][1]  ( .D(n496), .CLK(clk), .RSTB(n2334), .Q(reg15[1])
         );
  DFFARX1 \regf_reg[14][0]  ( .D(n495), .CLK(clk), .RSTB(n2334), .Q(reg15[0])
         );
  DFFARX1 \regf_reg[13][31]  ( .D(n494), .CLK(clk), .RSTB(n2334), .Q(reg14[31]) );
  DFFARX1 \regf_reg[13][30]  ( .D(n493), .CLK(clk), .RSTB(n2334), .Q(reg14[30]) );
  DFFARX1 \regf_reg[13][29]  ( .D(n492), .CLK(clk), .RSTB(n2334), .Q(reg14[29]) );
  DFFARX1 \regf_reg[13][28]  ( .D(n491), .CLK(clk), .RSTB(n2334), .Q(reg14[28]) );
  DFFARX1 \regf_reg[13][27]  ( .D(n490), .CLK(clk), .RSTB(n2334), .Q(reg14[27]) );
  DFFARX1 \regf_reg[13][26]  ( .D(n489), .CLK(clk), .RSTB(n2334), .Q(reg14[26]) );
  DFFARX1 \regf_reg[13][25]  ( .D(n488), .CLK(clk), .RSTB(n2334), .Q(reg14[25]) );
  DFFARX1 \regf_reg[13][24]  ( .D(n487), .CLK(clk), .RSTB(n2334), .Q(reg14[24]) );
  DFFARX1 \regf_reg[13][23]  ( .D(n486), .CLK(clk), .RSTB(n2333), .Q(reg14[23]) );
  DFFARX1 \regf_reg[13][22]  ( .D(n485), .CLK(clk), .RSTB(n2333), .Q(reg14[22]) );
  DFFARX1 \regf_reg[13][21]  ( .D(n484), .CLK(clk), .RSTB(n2333), .Q(reg14[21]) );
  DFFARX1 \regf_reg[13][20]  ( .D(n483), .CLK(clk), .RSTB(n2333), .Q(reg14[20]) );
  DFFARX1 \regf_reg[13][19]  ( .D(n482), .CLK(clk), .RSTB(n2333), .Q(reg14[19]) );
  DFFARX1 \regf_reg[13][18]  ( .D(n481), .CLK(clk), .RSTB(n2333), .Q(reg14[18]) );
  DFFARX1 \regf_reg[13][17]  ( .D(n480), .CLK(clk), .RSTB(n2333), .Q(reg14[17]) );
  DFFARX1 \regf_reg[13][16]  ( .D(n479), .CLK(clk), .RSTB(n2333), .Q(reg14[16]) );
  DFFARX1 \regf_reg[13][15]  ( .D(n478), .CLK(clk), .RSTB(n2333), .Q(reg14[15]) );
  DFFARX1 \regf_reg[13][14]  ( .D(n477), .CLK(clk), .RSTB(n2333), .Q(reg14[14]) );
  DFFARX1 \regf_reg[13][13]  ( .D(n476), .CLK(clk), .RSTB(n2333), .Q(reg14[13]) );
  DFFARX1 \regf_reg[13][12]  ( .D(n475), .CLK(clk), .RSTB(n2333), .Q(reg14[12]) );
  DFFARX1 \regf_reg[13][11]  ( .D(n474), .CLK(clk), .RSTB(n2332), .Q(reg14[11]) );
  DFFARX1 \regf_reg[13][10]  ( .D(n473), .CLK(clk), .RSTB(n2332), .Q(reg14[10]) );
  DFFARX1 \regf_reg[13][9]  ( .D(n472), .CLK(clk), .RSTB(n2332), .Q(reg14[9])
         );
  DFFARX1 \regf_reg[13][8]  ( .D(n471), .CLK(clk), .RSTB(n2332), .Q(reg14[8])
         );
  DFFARX1 \regf_reg[13][7]  ( .D(n470), .CLK(clk), .RSTB(n2332), .Q(reg14[7])
         );
  DFFARX1 \regf_reg[13][6]  ( .D(n469), .CLK(clk), .RSTB(n2332), .Q(reg14[6])
         );
  DFFARX1 \regf_reg[13][5]  ( .D(n468), .CLK(clk), .RSTB(n2332), .Q(reg14[5])
         );
  DFFARX1 \regf_reg[13][4]  ( .D(n467), .CLK(clk), .RSTB(n2332), .Q(reg14[4])
         );
  DFFARX1 \regf_reg[13][3]  ( .D(n466), .CLK(clk), .RSTB(n2332), .Q(reg14[3])
         );
  DFFARX1 \regf_reg[13][2]  ( .D(n465), .CLK(clk), .RSTB(n2332), .Q(reg14[2])
         );
  DFFARX1 \regf_reg[13][1]  ( .D(n464), .CLK(clk), .RSTB(n2332), .Q(reg14[1])
         );
  DFFARX1 \regf_reg[13][0]  ( .D(n463), .CLK(clk), .RSTB(n2332), .Q(reg14[0])
         );
  DFFARX1 \regf_reg[12][31]  ( .D(n462), .CLK(clk), .RSTB(n2331), .Q(reg13[31]) );
  DFFARX1 \regf_reg[12][30]  ( .D(n461), .CLK(clk), .RSTB(n2331), .Q(reg13[30]) );
  DFFARX1 \regf_reg[12][29]  ( .D(n460), .CLK(clk), .RSTB(n2331), .Q(reg13[29]) );
  DFFARX1 \regf_reg[12][28]  ( .D(n459), .CLK(clk), .RSTB(n2331), .Q(reg13[28]) );
  DFFARX1 \regf_reg[12][27]  ( .D(n458), .CLK(clk), .RSTB(n2331), .Q(reg13[27]) );
  DFFARX1 \regf_reg[12][26]  ( .D(n457), .CLK(clk), .RSTB(n2331), .Q(reg13[26]) );
  DFFARX1 \regf_reg[12][25]  ( .D(n456), .CLK(clk), .RSTB(n2331), .Q(reg13[25]) );
  DFFARX1 \regf_reg[12][24]  ( .D(n455), .CLK(clk), .RSTB(n2331), .Q(reg13[24]) );
  DFFARX1 \regf_reg[12][23]  ( .D(n454), .CLK(clk), .RSTB(n2331), .Q(reg13[23]) );
  DFFARX1 \regf_reg[12][22]  ( .D(n453), .CLK(clk), .RSTB(n2331), .Q(reg13[22]) );
  DFFARX1 \regf_reg[12][21]  ( .D(n452), .CLK(clk), .RSTB(n2331), .Q(reg13[21]) );
  DFFARX1 \regf_reg[12][20]  ( .D(n451), .CLK(clk), .RSTB(n2331), .Q(reg13[20]) );
  DFFARX1 \regf_reg[12][19]  ( .D(n450), .CLK(clk), .RSTB(n2330), .Q(reg13[19]) );
  DFFARX1 \regf_reg[12][18]  ( .D(n449), .CLK(clk), .RSTB(n2330), .Q(reg13[18]) );
  DFFARX1 \regf_reg[12][17]  ( .D(n448), .CLK(clk), .RSTB(n2330), .Q(reg13[17]) );
  DFFARX1 \regf_reg[12][16]  ( .D(n447), .CLK(clk), .RSTB(n2330), .Q(reg13[16]) );
  DFFARX1 \regf_reg[12][15]  ( .D(n446), .CLK(clk), .RSTB(n2330), .Q(reg13[15]) );
  DFFARX1 \regf_reg[12][14]  ( .D(n445), .CLK(clk), .RSTB(n2330), .Q(reg13[14]) );
  DFFARX1 \regf_reg[12][13]  ( .D(n444), .CLK(clk), .RSTB(n2330), .Q(reg13[13]) );
  DFFARX1 \regf_reg[12][12]  ( .D(n443), .CLK(clk), .RSTB(n2330), .Q(reg13[12]) );
  DFFARX1 \regf_reg[12][11]  ( .D(n442), .CLK(clk), .RSTB(n2330), .Q(reg13[11]) );
  DFFARX1 \regf_reg[12][10]  ( .D(n441), .CLK(clk), .RSTB(n2330), .Q(reg13[10]) );
  DFFARX1 \regf_reg[12][9]  ( .D(n440), .CLK(clk), .RSTB(n2330), .Q(reg13[9])
         );
  DFFARX1 \regf_reg[12][8]  ( .D(n439), .CLK(clk), .RSTB(n2330), .Q(reg13[8])
         );
  DFFARX1 \regf_reg[12][7]  ( .D(n438), .CLK(clk), .RSTB(n2329), .Q(reg13[7])
         );
  DFFARX1 \regf_reg[12][6]  ( .D(n437), .CLK(clk), .RSTB(n2329), .Q(reg13[6])
         );
  DFFARX1 \regf_reg[12][5]  ( .D(n436), .CLK(clk), .RSTB(n2329), .Q(reg13[5])
         );
  DFFARX1 \regf_reg[12][4]  ( .D(n435), .CLK(clk), .RSTB(n2329), .Q(reg13[4])
         );
  DFFARX1 \regf_reg[12][3]  ( .D(n434), .CLK(clk), .RSTB(n2329), .Q(reg13[3])
         );
  DFFARX1 \regf_reg[12][2]  ( .D(n433), .CLK(clk), .RSTB(n2329), .Q(reg13[2])
         );
  DFFARX1 \regf_reg[12][1]  ( .D(n432), .CLK(clk), .RSTB(n2329), .Q(reg13[1])
         );
  DFFARX1 \regf_reg[12][0]  ( .D(n431), .CLK(clk), .RSTB(n2329), .Q(reg13[0])
         );
  DFFARX1 \regf_reg[11][31]  ( .D(n430), .CLK(clk), .RSTB(n2329), .Q(reg12[31]) );
  DFFARX1 \regf_reg[11][30]  ( .D(n429), .CLK(clk), .RSTB(n2329), .Q(reg12[30]) );
  DFFARX1 \regf_reg[11][29]  ( .D(n428), .CLK(clk), .RSTB(n2329), .Q(reg12[29]) );
  DFFARX1 \regf_reg[11][28]  ( .D(n427), .CLK(clk), .RSTB(n2329), .Q(reg12[28]) );
  DFFARX1 \regf_reg[11][27]  ( .D(n426), .CLK(clk), .RSTB(n2328), .Q(reg12[27]) );
  DFFARX1 \regf_reg[11][26]  ( .D(n425), .CLK(clk), .RSTB(n2328), .Q(reg12[26]) );
  DFFARX1 \regf_reg[11][25]  ( .D(n424), .CLK(clk), .RSTB(n2328), .Q(reg12[25]) );
  DFFARX1 \regf_reg[11][24]  ( .D(n423), .CLK(clk), .RSTB(n2328), .Q(reg12[24]) );
  DFFARX1 \regf_reg[11][23]  ( .D(n422), .CLK(clk), .RSTB(n2328), .Q(reg12[23]) );
  DFFARX1 \regf_reg[11][22]  ( .D(n421), .CLK(clk), .RSTB(n2328), .Q(reg12[22]) );
  DFFARX1 \regf_reg[11][21]  ( .D(n420), .CLK(clk), .RSTB(n2328), .Q(reg12[21]) );
  DFFARX1 \regf_reg[11][20]  ( .D(n419), .CLK(clk), .RSTB(n2328), .Q(reg12[20]) );
  DFFARX1 \regf_reg[11][19]  ( .D(n418), .CLK(clk), .RSTB(n2328), .Q(reg12[19]) );
  DFFARX1 \regf_reg[11][18]  ( .D(n417), .CLK(clk), .RSTB(n2328), .Q(reg12[18]) );
  DFFARX1 \regf_reg[11][17]  ( .D(n416), .CLK(clk), .RSTB(n2328), .Q(reg12[17]) );
  DFFARX1 \regf_reg[11][16]  ( .D(n415), .CLK(clk), .RSTB(n2328), .Q(reg12[16]) );
  DFFARX1 \regf_reg[11][15]  ( .D(n414), .CLK(clk), .RSTB(n2327), .Q(reg12[15]) );
  DFFARX1 \regf_reg[11][14]  ( .D(n413), .CLK(clk), .RSTB(n2327), .Q(reg12[14]) );
  DFFARX1 \regf_reg[11][13]  ( .D(n412), .CLK(clk), .RSTB(n2327), .Q(reg12[13]) );
  DFFARX1 \regf_reg[11][12]  ( .D(n411), .CLK(clk), .RSTB(n2327), .Q(reg12[12]) );
  DFFARX1 \regf_reg[11][11]  ( .D(n410), .CLK(clk), .RSTB(n2327), .Q(reg12[11]) );
  DFFARX1 \regf_reg[11][10]  ( .D(n409), .CLK(clk), .RSTB(n2327), .Q(reg12[10]) );
  DFFARX1 \regf_reg[11][9]  ( .D(n408), .CLK(clk), .RSTB(n2327), .Q(reg12[9])
         );
  DFFARX1 \regf_reg[11][8]  ( .D(n407), .CLK(clk), .RSTB(n2327), .Q(reg12[8])
         );
  DFFARX1 \regf_reg[11][7]  ( .D(n406), .CLK(clk), .RSTB(n2327), .Q(reg12[7])
         );
  DFFARX1 \regf_reg[11][6]  ( .D(n405), .CLK(clk), .RSTB(n2327), .Q(reg12[6])
         );
  DFFARX1 \regf_reg[11][5]  ( .D(n404), .CLK(clk), .RSTB(n2327), .Q(reg12[5])
         );
  DFFARX1 \regf_reg[11][4]  ( .D(n403), .CLK(clk), .RSTB(n2327), .Q(reg12[4])
         );
  DFFARX1 \regf_reg[11][3]  ( .D(n402), .CLK(clk), .RSTB(n2326), .Q(reg12[3])
         );
  DFFARX1 \regf_reg[11][2]  ( .D(n401), .CLK(clk), .RSTB(n2326), .Q(reg12[2])
         );
  DFFARX1 \regf_reg[11][1]  ( .D(n400), .CLK(clk), .RSTB(n2326), .Q(reg12[1])
         );
  DFFARX1 \regf_reg[11][0]  ( .D(n399), .CLK(clk), .RSTB(n2326), .Q(reg12[0])
         );
  DFFARX1 \regf_reg[10][31]  ( .D(n398), .CLK(clk), .RSTB(n2326), .Q(reg11[31]) );
  DFFARX1 \regf_reg[10][30]  ( .D(n397), .CLK(clk), .RSTB(n2326), .Q(reg11[30]) );
  DFFARX1 \regf_reg[10][29]  ( .D(n396), .CLK(clk), .RSTB(n2326), .Q(reg11[29]) );
  DFFARX1 \regf_reg[10][28]  ( .D(n395), .CLK(clk), .RSTB(n2326), .Q(reg11[28]) );
  DFFARX1 \regf_reg[10][27]  ( .D(n394), .CLK(clk), .RSTB(n2326), .Q(reg11[27]) );
  DFFARX1 \regf_reg[10][26]  ( .D(n393), .CLK(clk), .RSTB(n2326), .Q(reg11[26]) );
  DFFARX1 \regf_reg[10][25]  ( .D(n392), .CLK(clk), .RSTB(n2326), .Q(reg11[25]) );
  DFFARX1 \regf_reg[10][24]  ( .D(n391), .CLK(clk), .RSTB(n2326), .Q(reg11[24]) );
  DFFARX1 \regf_reg[10][23]  ( .D(n390), .CLK(clk), .RSTB(n2325), .Q(reg11[23]) );
  DFFARX1 \regf_reg[10][22]  ( .D(n389), .CLK(clk), .RSTB(n2325), .Q(reg11[22]) );
  DFFARX1 \regf_reg[10][21]  ( .D(n388), .CLK(clk), .RSTB(n2325), .Q(reg11[21]) );
  DFFARX1 \regf_reg[10][20]  ( .D(n387), .CLK(clk), .RSTB(n2325), .Q(reg11[20]) );
  DFFARX1 \regf_reg[10][19]  ( .D(n386), .CLK(clk), .RSTB(n2325), .Q(reg11[19]) );
  DFFARX1 \regf_reg[10][18]  ( .D(n385), .CLK(clk), .RSTB(n2325), .Q(reg11[18]) );
  DFFARX1 \regf_reg[10][17]  ( .D(n384), .CLK(clk), .RSTB(n2325), .Q(reg11[17]) );
  DFFARX1 \regf_reg[10][16]  ( .D(n383), .CLK(clk), .RSTB(n2325), .Q(reg11[16]) );
  DFFARX1 \regf_reg[10][15]  ( .D(n382), .CLK(clk), .RSTB(n2325), .Q(reg11[15]) );
  DFFARX1 \regf_reg[10][14]  ( .D(n381), .CLK(clk), .RSTB(n2325), .Q(reg11[14]) );
  DFFARX1 \regf_reg[10][13]  ( .D(n380), .CLK(clk), .RSTB(n2325), .Q(reg11[13]) );
  DFFARX1 \regf_reg[10][12]  ( .D(n379), .CLK(clk), .RSTB(n2325), .Q(reg11[12]) );
  DFFARX1 \regf_reg[10][11]  ( .D(n378), .CLK(clk), .RSTB(n2324), .Q(reg11[11]) );
  DFFARX1 \regf_reg[10][10]  ( .D(n377), .CLK(clk), .RSTB(n2324), .Q(reg11[10]) );
  DFFARX1 \regf_reg[10][9]  ( .D(n376), .CLK(clk), .RSTB(n2324), .Q(reg11[9])
         );
  DFFARX1 \regf_reg[10][8]  ( .D(n375), .CLK(clk), .RSTB(n2324), .Q(reg11[8])
         );
  DFFARX1 \regf_reg[10][7]  ( .D(n374), .CLK(clk), .RSTB(n2324), .Q(reg11[7])
         );
  DFFARX1 \regf_reg[10][6]  ( .D(n373), .CLK(clk), .RSTB(n2324), .Q(reg11[6])
         );
  DFFARX1 \regf_reg[10][5]  ( .D(n372), .CLK(clk), .RSTB(n2324), .Q(reg11[5])
         );
  DFFARX1 \regf_reg[10][4]  ( .D(n371), .CLK(clk), .RSTB(n2324), .Q(reg11[4])
         );
  DFFARX1 \regf_reg[10][3]  ( .D(n370), .CLK(clk), .RSTB(n2324), .Q(reg11[3])
         );
  DFFARX1 \regf_reg[10][2]  ( .D(n369), .CLK(clk), .RSTB(n2324), .Q(reg11[2])
         );
  DFFARX1 \regf_reg[10][1]  ( .D(n368), .CLK(clk), .RSTB(n2324), .Q(reg11[1])
         );
  DFFARX1 \regf_reg[10][0]  ( .D(n367), .CLK(clk), .RSTB(n2324), .Q(reg11[0])
         );
  DFFARX1 \regf_reg[9][31]  ( .D(n366), .CLK(clk), .RSTB(n2323), .Q(reg10[31])
         );
  DFFARX1 \regf_reg[9][30]  ( .D(n365), .CLK(clk), .RSTB(n2323), .Q(reg10[30])
         );
  DFFARX1 \regf_reg[9][29]  ( .D(n364), .CLK(clk), .RSTB(n2323), .Q(reg10[29])
         );
  DFFARX1 \regf_reg[9][28]  ( .D(n363), .CLK(clk), .RSTB(n2323), .Q(reg10[28])
         );
  DFFARX1 \regf_reg[9][27]  ( .D(n362), .CLK(clk), .RSTB(n2323), .Q(reg10[27])
         );
  DFFARX1 \regf_reg[9][26]  ( .D(n361), .CLK(clk), .RSTB(n2323), .Q(reg10[26])
         );
  DFFARX1 \regf_reg[9][25]  ( .D(n360), .CLK(clk), .RSTB(n2323), .Q(reg10[25])
         );
  DFFARX1 \regf_reg[9][24]  ( .D(n359), .CLK(clk), .RSTB(n2323), .Q(reg10[24])
         );
  DFFARX1 \regf_reg[9][23]  ( .D(n358), .CLK(clk), .RSTB(n2323), .Q(reg10[23])
         );
  DFFARX1 \regf_reg[9][22]  ( .D(n357), .CLK(clk), .RSTB(n2323), .Q(reg10[22])
         );
  DFFARX1 \regf_reg[9][21]  ( .D(n356), .CLK(clk), .RSTB(n2323), .Q(reg10[21])
         );
  DFFARX1 \regf_reg[9][20]  ( .D(n355), .CLK(clk), .RSTB(n2323), .Q(reg10[20])
         );
  DFFARX1 \regf_reg[9][19]  ( .D(n354), .CLK(clk), .RSTB(n2322), .Q(reg10[19])
         );
  DFFARX1 \regf_reg[9][18]  ( .D(n353), .CLK(clk), .RSTB(n2322), .Q(reg10[18])
         );
  DFFARX1 \regf_reg[9][17]  ( .D(n352), .CLK(clk), .RSTB(n2322), .Q(reg10[17])
         );
  DFFARX1 \regf_reg[9][16]  ( .D(n351), .CLK(clk), .RSTB(n2322), .Q(reg10[16])
         );
  DFFARX1 \regf_reg[9][15]  ( .D(n350), .CLK(clk), .RSTB(n2322), .Q(reg10[15])
         );
  DFFARX1 \regf_reg[9][14]  ( .D(n349), .CLK(clk), .RSTB(n2322), .Q(reg10[14])
         );
  DFFARX1 \regf_reg[9][13]  ( .D(n348), .CLK(clk), .RSTB(n2322), .Q(reg10[13])
         );
  DFFARX1 \regf_reg[9][12]  ( .D(n347), .CLK(clk), .RSTB(n2322), .Q(reg10[12])
         );
  DFFARX1 \regf_reg[9][11]  ( .D(n346), .CLK(clk), .RSTB(n2322), .Q(reg10[11])
         );
  DFFARX1 \regf_reg[9][10]  ( .D(n345), .CLK(clk), .RSTB(n2322), .Q(reg10[10])
         );
  DFFARX1 \regf_reg[9][9]  ( .D(n344), .CLK(clk), .RSTB(n2322), .Q(reg10[9])
         );
  DFFARX1 \regf_reg[9][8]  ( .D(n343), .CLK(clk), .RSTB(n2322), .Q(reg10[8])
         );
  DFFARX1 \regf_reg[9][7]  ( .D(n342), .CLK(clk), .RSTB(n2321), .Q(reg10[7])
         );
  DFFARX1 \regf_reg[9][6]  ( .D(n341), .CLK(clk), .RSTB(n2321), .Q(reg10[6])
         );
  DFFARX1 \regf_reg[9][5]  ( .D(n340), .CLK(clk), .RSTB(n2321), .Q(reg10[5])
         );
  DFFARX1 \regf_reg[9][4]  ( .D(n339), .CLK(clk), .RSTB(n2321), .Q(reg10[4])
         );
  DFFARX1 \regf_reg[9][3]  ( .D(n338), .CLK(clk), .RSTB(n2321), .Q(reg10[3])
         );
  DFFARX1 \regf_reg[9][2]  ( .D(n337), .CLK(clk), .RSTB(n2321), .Q(reg10[2])
         );
  DFFARX1 \regf_reg[9][1]  ( .D(n336), .CLK(clk), .RSTB(n2321), .Q(reg10[1])
         );
  DFFARX1 \regf_reg[9][0]  ( .D(n335), .CLK(clk), .RSTB(n2321), .Q(reg10[0])
         );
  DFFARX1 \regf_reg[8][31]  ( .D(n334), .CLK(clk), .RSTB(n2321), .Q(reg9[31])
         );
  DFFARX1 \regf_reg[8][30]  ( .D(n333), .CLK(clk), .RSTB(n2321), .Q(reg9[30])
         );
  DFFARX1 \regf_reg[8][29]  ( .D(n332), .CLK(clk), .RSTB(n2321), .Q(reg9[29])
         );
  DFFARX1 \regf_reg[8][28]  ( .D(n331), .CLK(clk), .RSTB(n2321), .Q(reg9[28])
         );
  DFFARX1 \regf_reg[8][27]  ( .D(n330), .CLK(clk), .RSTB(n2320), .Q(reg9[27])
         );
  DFFARX1 \regf_reg[8][26]  ( .D(n329), .CLK(clk), .RSTB(n2320), .Q(reg9[26])
         );
  DFFARX1 \regf_reg[8][25]  ( .D(n328), .CLK(clk), .RSTB(n2320), .Q(reg9[25])
         );
  DFFARX1 \regf_reg[8][24]  ( .D(n327), .CLK(clk), .RSTB(n2320), .Q(reg9[24])
         );
  DFFARX1 \regf_reg[8][23]  ( .D(n326), .CLK(clk), .RSTB(n2320), .Q(reg9[23])
         );
  DFFARX1 \regf_reg[8][22]  ( .D(n325), .CLK(clk), .RSTB(n2320), .Q(reg9[22])
         );
  DFFARX1 \regf_reg[8][21]  ( .D(n324), .CLK(clk), .RSTB(n2320), .Q(reg9[21])
         );
  DFFARX1 \regf_reg[8][20]  ( .D(n323), .CLK(clk), .RSTB(n2320), .Q(reg9[20])
         );
  DFFARX1 \regf_reg[8][19]  ( .D(n322), .CLK(clk), .RSTB(n2320), .Q(reg9[19])
         );
  DFFARX1 \regf_reg[8][18]  ( .D(n321), .CLK(clk), .RSTB(n2320), .Q(reg9[18])
         );
  DFFARX1 \regf_reg[8][17]  ( .D(n320), .CLK(clk), .RSTB(n2320), .Q(reg9[17])
         );
  DFFARX1 \regf_reg[8][16]  ( .D(n319), .CLK(clk), .RSTB(n2320), .Q(reg9[16])
         );
  DFFARX1 \regf_reg[8][15]  ( .D(n318), .CLK(clk), .RSTB(n2319), .Q(reg9[15])
         );
  DFFARX1 \regf_reg[8][14]  ( .D(n317), .CLK(clk), .RSTB(n2319), .Q(reg9[14])
         );
  DFFARX1 \regf_reg[8][13]  ( .D(n316), .CLK(clk), .RSTB(n2319), .Q(reg9[13])
         );
  DFFARX1 \regf_reg[8][12]  ( .D(n315), .CLK(clk), .RSTB(n2319), .Q(reg9[12])
         );
  DFFARX1 \regf_reg[8][11]  ( .D(n314), .CLK(clk), .RSTB(n2319), .Q(reg9[11])
         );
  DFFARX1 \regf_reg[8][10]  ( .D(n313), .CLK(clk), .RSTB(n2319), .Q(reg9[10])
         );
  DFFARX1 \regf_reg[8][9]  ( .D(n312), .CLK(clk), .RSTB(n2319), .Q(reg9[9]) );
  DFFARX1 \regf_reg[8][8]  ( .D(n311), .CLK(clk), .RSTB(n2319), .Q(reg9[8]) );
  DFFARX1 \regf_reg[8][7]  ( .D(n310), .CLK(clk), .RSTB(n2319), .Q(reg9[7]) );
  DFFARX1 \regf_reg[8][6]  ( .D(n309), .CLK(clk), .RSTB(n2319), .Q(reg9[6]) );
  DFFARX1 \regf_reg[8][5]  ( .D(n308), .CLK(clk), .RSTB(n2319), .Q(reg9[5]) );
  DFFARX1 \regf_reg[8][4]  ( .D(n307), .CLK(clk), .RSTB(n2319), .Q(reg9[4]) );
  DFFARX1 \regf_reg[8][3]  ( .D(n306), .CLK(clk), .RSTB(n2318), .Q(reg9[3]) );
  DFFARX1 \regf_reg[8][2]  ( .D(n305), .CLK(clk), .RSTB(n2318), .Q(reg9[2]) );
  DFFARX1 \regf_reg[8][1]  ( .D(n304), .CLK(clk), .RSTB(n2318), .Q(reg9[1]) );
  DFFARX1 \regf_reg[8][0]  ( .D(n303), .CLK(clk), .RSTB(n2318), .Q(reg9[0]) );
  DFFARX1 \regf_reg[7][31]  ( .D(n302), .CLK(clk), .RSTB(n2318), .Q(reg8[31])
         );
  DFFARX1 \regf_reg[7][30]  ( .D(n301), .CLK(clk), .RSTB(n2318), .Q(reg8[30])
         );
  DFFARX1 \regf_reg[7][29]  ( .D(n300), .CLK(clk), .RSTB(n2318), .Q(reg8[29])
         );
  DFFARX1 \regf_reg[7][28]  ( .D(n299), .CLK(clk), .RSTB(n2318), .Q(reg8[28])
         );
  DFFARX1 \regf_reg[7][27]  ( .D(n298), .CLK(clk), .RSTB(n2318), .Q(reg8[27])
         );
  DFFARX1 \regf_reg[7][26]  ( .D(n297), .CLK(clk), .RSTB(n2318), .Q(reg8[26])
         );
  DFFARX1 \regf_reg[7][25]  ( .D(n296), .CLK(clk), .RSTB(n2318), .Q(reg8[25])
         );
  DFFARX1 \regf_reg[7][24]  ( .D(n295), .CLK(clk), .RSTB(n2318), .Q(reg8[24])
         );
  DFFARX1 \regf_reg[7][23]  ( .D(n294), .CLK(clk), .RSTB(n2317), .Q(reg8[23])
         );
  DFFARX1 \regf_reg[7][22]  ( .D(n293), .CLK(clk), .RSTB(n2317), .Q(reg8[22])
         );
  DFFARX1 \regf_reg[7][21]  ( .D(n292), .CLK(clk), .RSTB(n2317), .Q(reg8[21])
         );
  DFFARX1 \regf_reg[7][20]  ( .D(n291), .CLK(clk), .RSTB(n2317), .Q(reg8[20])
         );
  DFFARX1 \regf_reg[7][19]  ( .D(n290), .CLK(clk), .RSTB(n2317), .Q(reg8[19])
         );
  DFFARX1 \regf_reg[7][18]  ( .D(n289), .CLK(clk), .RSTB(n2317), .Q(reg8[18])
         );
  DFFARX1 \regf_reg[7][17]  ( .D(n288), .CLK(clk), .RSTB(n2317), .Q(reg8[17])
         );
  DFFARX1 \regf_reg[7][16]  ( .D(n287), .CLK(clk), .RSTB(n2317), .Q(reg8[16])
         );
  DFFARX1 \regf_reg[7][15]  ( .D(n286), .CLK(clk), .RSTB(n2317), .Q(reg8[15])
         );
  DFFARX1 \regf_reg[7][14]  ( .D(n285), .CLK(clk), .RSTB(n2317), .Q(reg8[14])
         );
  DFFARX1 \regf_reg[7][13]  ( .D(n284), .CLK(clk), .RSTB(n2317), .Q(reg8[13])
         );
  DFFARX1 \regf_reg[7][12]  ( .D(n283), .CLK(clk), .RSTB(n2317), .Q(reg8[12])
         );
  DFFARX1 \regf_reg[7][11]  ( .D(n282), .CLK(clk), .RSTB(n2316), .Q(reg8[11])
         );
  DFFARX1 \regf_reg[7][10]  ( .D(n281), .CLK(clk), .RSTB(n2316), .Q(reg8[10])
         );
  DFFARX1 \regf_reg[7][9]  ( .D(n280), .CLK(clk), .RSTB(n2316), .Q(reg8[9]) );
  DFFARX1 \regf_reg[7][8]  ( .D(n279), .CLK(clk), .RSTB(n2316), .Q(reg8[8]) );
  DFFARX1 \regf_reg[7][7]  ( .D(n278), .CLK(clk), .RSTB(n2316), .Q(reg8[7]) );
  DFFARX1 \regf_reg[7][6]  ( .D(n277), .CLK(clk), .RSTB(n2316), .Q(reg8[6]) );
  DFFARX1 \regf_reg[7][5]  ( .D(n276), .CLK(clk), .RSTB(n2316), .Q(reg8[5]) );
  DFFARX1 \regf_reg[7][4]  ( .D(n275), .CLK(clk), .RSTB(n2316), .Q(reg8[4]) );
  DFFARX1 \regf_reg[7][3]  ( .D(n274), .CLK(clk), .RSTB(n2316), .Q(reg8[3]) );
  DFFARX1 \regf_reg[7][2]  ( .D(n273), .CLK(clk), .RSTB(n2316), .Q(reg8[2]) );
  DFFARX1 \regf_reg[7][1]  ( .D(n272), .CLK(clk), .RSTB(n2316), .Q(reg8[1]) );
  DFFARX1 \regf_reg[7][0]  ( .D(n271), .CLK(clk), .RSTB(n2316), .Q(reg8[0]) );
  DFFARX1 \regf_reg[6][31]  ( .D(n270), .CLK(clk), .RSTB(n2315), .Q(reg7[31])
         );
  DFFARX1 \regf_reg[6][30]  ( .D(n269), .CLK(clk), .RSTB(n2315), .Q(reg7[30])
         );
  DFFARX1 \regf_reg[6][29]  ( .D(n268), .CLK(clk), .RSTB(n2315), .Q(reg7[29])
         );
  DFFARX1 \regf_reg[6][28]  ( .D(n267), .CLK(clk), .RSTB(n2315), .Q(reg7[28])
         );
  DFFARX1 \regf_reg[6][27]  ( .D(n266), .CLK(clk), .RSTB(n2315), .Q(reg7[27])
         );
  DFFARX1 \regf_reg[6][26]  ( .D(n265), .CLK(clk), .RSTB(n2315), .Q(reg7[26])
         );
  DFFARX1 \regf_reg[6][25]  ( .D(n264), .CLK(clk), .RSTB(n2315), .Q(reg7[25])
         );
  DFFARX1 \regf_reg[6][24]  ( .D(n263), .CLK(clk), .RSTB(n2315), .Q(reg7[24])
         );
  DFFARX1 \regf_reg[6][23]  ( .D(n262), .CLK(clk), .RSTB(n2315), .Q(reg7[23])
         );
  DFFARX1 \regf_reg[6][22]  ( .D(n261), .CLK(clk), .RSTB(n2315), .Q(reg7[22])
         );
  DFFARX1 \regf_reg[6][21]  ( .D(n260), .CLK(clk), .RSTB(n2315), .Q(reg7[21])
         );
  DFFARX1 \regf_reg[6][20]  ( .D(n259), .CLK(clk), .RSTB(n2315), .Q(reg7[20])
         );
  DFFARX1 \regf_reg[6][19]  ( .D(n258), .CLK(clk), .RSTB(n2314), .Q(reg7[19])
         );
  DFFARX1 \regf_reg[6][18]  ( .D(n257), .CLK(clk), .RSTB(n2314), .Q(reg7[18])
         );
  DFFARX1 \regf_reg[6][17]  ( .D(n256), .CLK(clk), .RSTB(n2314), .Q(reg7[17])
         );
  DFFARX1 \regf_reg[6][16]  ( .D(n255), .CLK(clk), .RSTB(n2314), .Q(reg7[16])
         );
  DFFARX1 \regf_reg[6][15]  ( .D(n254), .CLK(clk), .RSTB(n2314), .Q(reg7[15])
         );
  DFFARX1 \regf_reg[6][14]  ( .D(n253), .CLK(clk), .RSTB(n2314), .Q(reg7[14])
         );
  DFFARX1 \regf_reg[6][13]  ( .D(n252), .CLK(clk), .RSTB(n2314), .Q(reg7[13])
         );
  DFFARX1 \regf_reg[6][12]  ( .D(n251), .CLK(clk), .RSTB(n2314), .Q(reg7[12])
         );
  DFFARX1 \regf_reg[6][11]  ( .D(n250), .CLK(clk), .RSTB(n2314), .Q(reg7[11])
         );
  DFFARX1 \regf_reg[6][10]  ( .D(n249), .CLK(clk), .RSTB(n2314), .Q(reg7[10])
         );
  DFFARX1 \regf_reg[6][9]  ( .D(n248), .CLK(clk), .RSTB(n2314), .Q(reg7[9]) );
  DFFARX1 \regf_reg[6][8]  ( .D(n247), .CLK(clk), .RSTB(n2314), .Q(reg7[8]) );
  DFFARX1 \regf_reg[6][7]  ( .D(n246), .CLK(clk), .RSTB(n2313), .Q(reg7[7]) );
  DFFARX1 \regf_reg[6][6]  ( .D(n245), .CLK(clk), .RSTB(n2313), .Q(reg7[6]) );
  DFFARX1 \regf_reg[6][5]  ( .D(n244), .CLK(clk), .RSTB(n2313), .Q(reg7[5]) );
  DFFARX1 \regf_reg[6][4]  ( .D(n243), .CLK(clk), .RSTB(n2313), .Q(reg7[4]) );
  DFFARX1 \regf_reg[6][3]  ( .D(n242), .CLK(clk), .RSTB(n2313), .Q(reg7[3]) );
  DFFARX1 \regf_reg[6][2]  ( .D(n241), .CLK(clk), .RSTB(n2313), .Q(reg7[2]) );
  DFFARX1 \regf_reg[6][1]  ( .D(n240), .CLK(clk), .RSTB(n2313), .Q(reg7[1]) );
  DFFARX1 \regf_reg[6][0]  ( .D(n239), .CLK(clk), .RSTB(n2313), .Q(reg7[0]) );
  DFFARX1 \regf_reg[5][31]  ( .D(n238), .CLK(clk), .RSTB(n2313), .Q(reg6[31])
         );
  DFFARX1 \regf_reg[5][30]  ( .D(n237), .CLK(clk), .RSTB(n2313), .Q(reg6[30])
         );
  DFFARX1 \regf_reg[5][29]  ( .D(n236), .CLK(clk), .RSTB(n2313), .Q(reg6[29])
         );
  DFFARX1 \regf_reg[5][28]  ( .D(n235), .CLK(clk), .RSTB(n2313), .Q(reg6[28])
         );
  DFFARX1 \regf_reg[5][27]  ( .D(n234), .CLK(clk), .RSTB(n2312), .Q(reg6[27])
         );
  DFFARX1 \regf_reg[5][26]  ( .D(n233), .CLK(clk), .RSTB(n2312), .Q(reg6[26])
         );
  DFFARX1 \regf_reg[5][25]  ( .D(n232), .CLK(clk), .RSTB(n2312), .Q(reg6[25])
         );
  DFFARX1 \regf_reg[5][24]  ( .D(n231), .CLK(clk), .RSTB(n2312), .Q(reg6[24])
         );
  DFFARX1 \regf_reg[5][23]  ( .D(n230), .CLK(clk), .RSTB(n2312), .Q(reg6[23])
         );
  DFFARX1 \regf_reg[5][22]  ( .D(n229), .CLK(clk), .RSTB(n2312), .Q(reg6[22])
         );
  DFFARX1 \regf_reg[5][21]  ( .D(n228), .CLK(clk), .RSTB(n2312), .Q(reg6[21])
         );
  DFFARX1 \regf_reg[5][20]  ( .D(n227), .CLK(clk), .RSTB(n2312), .Q(reg6[20])
         );
  DFFARX1 \regf_reg[5][19]  ( .D(n226), .CLK(clk), .RSTB(n2312), .Q(reg6[19])
         );
  DFFARX1 \regf_reg[5][18]  ( .D(n225), .CLK(clk), .RSTB(n2312), .Q(reg6[18])
         );
  DFFARX1 \regf_reg[5][17]  ( .D(n224), .CLK(clk), .RSTB(n2312), .Q(reg6[17])
         );
  DFFARX1 \regf_reg[5][16]  ( .D(n223), .CLK(clk), .RSTB(n2312), .Q(reg6[16])
         );
  DFFARX1 \regf_reg[5][15]  ( .D(n222), .CLK(clk), .RSTB(n2311), .Q(reg6[15])
         );
  DFFARX1 \regf_reg[5][14]  ( .D(n221), .CLK(clk), .RSTB(n2311), .Q(reg6[14])
         );
  DFFARX1 \regf_reg[5][13]  ( .D(n220), .CLK(clk), .RSTB(n2311), .Q(reg6[13])
         );
  DFFARX1 \regf_reg[5][12]  ( .D(n219), .CLK(clk), .RSTB(n2311), .Q(reg6[12])
         );
  DFFARX1 \regf_reg[5][11]  ( .D(n218), .CLK(clk), .RSTB(n2311), .Q(reg6[11])
         );
  DFFARX1 \regf_reg[5][10]  ( .D(n217), .CLK(clk), .RSTB(n2311), .Q(reg6[10])
         );
  DFFARX1 \regf_reg[5][9]  ( .D(n216), .CLK(clk), .RSTB(n2311), .Q(reg6[9]) );
  DFFARX1 \regf_reg[5][8]  ( .D(n215), .CLK(clk), .RSTB(n2311), .Q(reg6[8]) );
  DFFARX1 \regf_reg[5][7]  ( .D(n214), .CLK(clk), .RSTB(n2311), .Q(reg6[7]) );
  DFFARX1 \regf_reg[5][6]  ( .D(n213), .CLK(clk), .RSTB(n2311), .Q(reg6[6]) );
  DFFARX1 \regf_reg[5][5]  ( .D(n212), .CLK(clk), .RSTB(n2311), .Q(reg6[5]) );
  DFFARX1 \regf_reg[5][4]  ( .D(n211), .CLK(clk), .RSTB(n2311), .Q(reg6[4]) );
  DFFARX1 \regf_reg[5][3]  ( .D(n210), .CLK(clk), .RSTB(n2310), .Q(reg6[3]) );
  DFFARX1 \regf_reg[5][2]  ( .D(n209), .CLK(clk), .RSTB(n2310), .Q(reg6[2]) );
  DFFARX1 \regf_reg[5][1]  ( .D(n208), .CLK(clk), .RSTB(n2310), .Q(reg6[1]) );
  DFFARX1 \regf_reg[5][0]  ( .D(n207), .CLK(clk), .RSTB(n2310), .Q(reg6[0]) );
  DFFARX1 \regf_reg[4][31]  ( .D(n206), .CLK(clk), .RSTB(n2310), .Q(reg5[31])
         );
  DFFARX1 \regf_reg[4][30]  ( .D(n205), .CLK(clk), .RSTB(n2310), .Q(reg5[30])
         );
  DFFARX1 \regf_reg[4][29]  ( .D(n204), .CLK(clk), .RSTB(n2310), .Q(reg5[29])
         );
  DFFARX1 \regf_reg[4][28]  ( .D(n203), .CLK(clk), .RSTB(n2310), .Q(reg5[28])
         );
  DFFARX1 \regf_reg[4][27]  ( .D(n202), .CLK(clk), .RSTB(n2310), .Q(reg5[27])
         );
  DFFARX1 \regf_reg[4][26]  ( .D(n201), .CLK(clk), .RSTB(n2310), .Q(reg5[26])
         );
  DFFARX1 \regf_reg[4][25]  ( .D(n200), .CLK(clk), .RSTB(n2310), .Q(reg5[25])
         );
  DFFARX1 \regf_reg[4][24]  ( .D(n199), .CLK(clk), .RSTB(n2310), .Q(reg5[24])
         );
  DFFARX1 \regf_reg[4][23]  ( .D(n198), .CLK(clk), .RSTB(n2309), .Q(reg5[23])
         );
  DFFARX1 \regf_reg[4][22]  ( .D(n197), .CLK(clk), .RSTB(n2309), .Q(reg5[22])
         );
  DFFARX1 \regf_reg[4][21]  ( .D(n196), .CLK(clk), .RSTB(n2309), .Q(reg5[21])
         );
  DFFARX1 \regf_reg[4][20]  ( .D(n195), .CLK(clk), .RSTB(n2309), .Q(reg5[20])
         );
  DFFARX1 \regf_reg[4][19]  ( .D(n194), .CLK(clk), .RSTB(n2309), .Q(reg5[19])
         );
  DFFARX1 \regf_reg[4][18]  ( .D(n193), .CLK(clk), .RSTB(n2309), .Q(reg5[18])
         );
  DFFARX1 \regf_reg[4][17]  ( .D(n192), .CLK(clk), .RSTB(n2309), .Q(reg5[17])
         );
  DFFARX1 \regf_reg[4][16]  ( .D(n191), .CLK(clk), .RSTB(n2309), .Q(reg5[16])
         );
  DFFARX1 \regf_reg[4][15]  ( .D(n190), .CLK(clk), .RSTB(n2309), .Q(reg5[15])
         );
  DFFARX1 \regf_reg[4][14]  ( .D(n189), .CLK(clk), .RSTB(n2309), .Q(reg5[14])
         );
  DFFARX1 \regf_reg[4][13]  ( .D(n188), .CLK(clk), .RSTB(n2309), .Q(reg5[13])
         );
  DFFARX1 \regf_reg[4][12]  ( .D(n187), .CLK(clk), .RSTB(n2309), .Q(reg5[12])
         );
  DFFARX1 \regf_reg[4][11]  ( .D(n186), .CLK(clk), .RSTB(n2308), .Q(reg5[11])
         );
  DFFARX1 \regf_reg[4][10]  ( .D(n185), .CLK(clk), .RSTB(n2308), .Q(reg5[10])
         );
  DFFARX1 \regf_reg[4][9]  ( .D(n184), .CLK(clk), .RSTB(n2308), .Q(reg5[9]) );
  DFFARX1 \regf_reg[4][8]  ( .D(n183), .CLK(clk), .RSTB(n2308), .Q(reg5[8]) );
  DFFARX1 \regf_reg[4][7]  ( .D(n182), .CLK(clk), .RSTB(n2308), .Q(reg5[7]) );
  DFFARX1 \regf_reg[4][6]  ( .D(n181), .CLK(clk), .RSTB(n2308), .Q(reg5[6]) );
  DFFARX1 \regf_reg[4][5]  ( .D(n180), .CLK(clk), .RSTB(n2308), .Q(reg5[5]) );
  DFFARX1 \regf_reg[4][4]  ( .D(n179), .CLK(clk), .RSTB(n2308), .Q(reg5[4]) );
  DFFARX1 \regf_reg[4][3]  ( .D(n178), .CLK(clk), .RSTB(n2308), .Q(reg5[3]) );
  DFFARX1 \regf_reg[4][2]  ( .D(n177), .CLK(clk), .RSTB(n2308), .Q(reg5[2]) );
  DFFARX1 \regf_reg[4][1]  ( .D(n176), .CLK(clk), .RSTB(n2308), .Q(reg5[1]) );
  DFFARX1 \regf_reg[4][0]  ( .D(n175), .CLK(clk), .RSTB(n2308), .Q(reg5[0]) );
  DFFARX1 \regf_reg[3][31]  ( .D(n174), .CLK(clk), .RSTB(n2307), .Q(reg4[31])
         );
  DFFARX1 \regf_reg[3][30]  ( .D(n173), .CLK(clk), .RSTB(n2307), .Q(reg4[30])
         );
  DFFARX1 \regf_reg[3][29]  ( .D(n172), .CLK(clk), .RSTB(n2307), .Q(reg4[29])
         );
  DFFARX1 \regf_reg[3][28]  ( .D(n171), .CLK(clk), .RSTB(n2307), .Q(reg4[28])
         );
  DFFARX1 \regf_reg[3][27]  ( .D(n170), .CLK(clk), .RSTB(n2307), .Q(reg4[27])
         );
  DFFARX1 \regf_reg[3][26]  ( .D(n169), .CLK(clk), .RSTB(n2307), .Q(reg4[26])
         );
  DFFARX1 \regf_reg[3][25]  ( .D(n168), .CLK(clk), .RSTB(n2307), .Q(reg4[25])
         );
  DFFARX1 \regf_reg[3][24]  ( .D(n167), .CLK(clk), .RSTB(n2307), .Q(reg4[24])
         );
  DFFARX1 \regf_reg[3][23]  ( .D(n166), .CLK(clk), .RSTB(n2307), .Q(reg4[23])
         );
  DFFARX1 \regf_reg[3][22]  ( .D(n165), .CLK(clk), .RSTB(n2307), .Q(reg4[22])
         );
  DFFARX1 \regf_reg[3][21]  ( .D(n164), .CLK(clk), .RSTB(n2307), .Q(reg4[21])
         );
  DFFARX1 \regf_reg[3][20]  ( .D(n163), .CLK(clk), .RSTB(n2307), .Q(reg4[20])
         );
  DFFARX1 \regf_reg[3][19]  ( .D(n162), .CLK(clk), .RSTB(n2306), .Q(reg4[19])
         );
  DFFARX1 \regf_reg[3][18]  ( .D(n161), .CLK(clk), .RSTB(n2306), .Q(reg4[18])
         );
  DFFARX1 \regf_reg[3][17]  ( .D(n160), .CLK(clk), .RSTB(n2306), .Q(reg4[17])
         );
  DFFARX1 \regf_reg[3][16]  ( .D(n159), .CLK(clk), .RSTB(n2306), .Q(reg4[16])
         );
  DFFARX1 \regf_reg[3][15]  ( .D(n158), .CLK(clk), .RSTB(n2306), .Q(reg4[15])
         );
  DFFARX1 \regf_reg[3][14]  ( .D(n157), .CLK(clk), .RSTB(n2306), .Q(reg4[14])
         );
  DFFARX1 \regf_reg[3][13]  ( .D(n156), .CLK(clk), .RSTB(n2306), .Q(reg4[13])
         );
  DFFARX1 \regf_reg[3][12]  ( .D(n155), .CLK(clk), .RSTB(n2306), .Q(reg4[12])
         );
  DFFARX1 \regf_reg[3][11]  ( .D(n154), .CLK(clk), .RSTB(n2306), .Q(reg4[11])
         );
  DFFARX1 \regf_reg[3][10]  ( .D(n153), .CLK(clk), .RSTB(n2306), .Q(reg4[10])
         );
  DFFARX1 \regf_reg[3][9]  ( .D(n152), .CLK(clk), .RSTB(n2306), .Q(reg4[9]) );
  DFFARX1 \regf_reg[3][8]  ( .D(n151), .CLK(clk), .RSTB(n2306), .Q(reg4[8]) );
  DFFARX1 \regf_reg[3][7]  ( .D(n150), .CLK(clk), .RSTB(n2305), .Q(reg4[7]) );
  DFFARX1 \regf_reg[3][6]  ( .D(n149), .CLK(clk), .RSTB(n2305), .Q(reg4[6]) );
  DFFARX1 \regf_reg[3][5]  ( .D(n148), .CLK(clk), .RSTB(n2305), .Q(reg4[5]) );
  DFFARX1 \regf_reg[3][4]  ( .D(n147), .CLK(clk), .RSTB(n2305), .Q(reg4[4]) );
  DFFARX1 \regf_reg[3][3]  ( .D(n146), .CLK(clk), .RSTB(n2305), .Q(reg4[3]) );
  DFFARX1 \regf_reg[3][2]  ( .D(n145), .CLK(clk), .RSTB(n2305), .Q(reg4[2]) );
  DFFARX1 \regf_reg[3][1]  ( .D(n144), .CLK(clk), .RSTB(n2305), .Q(reg4[1]) );
  DFFARX1 \regf_reg[3][0]  ( .D(n143), .CLK(clk), .RSTB(n2305), .Q(reg4[0]) );
  DFFARX1 \regf_reg[2][31]  ( .D(n142), .CLK(clk), .RSTB(n2305), .Q(reg3[31])
         );
  DFFARX1 \regf_reg[2][30]  ( .D(n141), .CLK(clk), .RSTB(n2305), .Q(reg3[30])
         );
  DFFARX1 \regf_reg[2][29]  ( .D(n140), .CLK(clk), .RSTB(n2305), .Q(reg3[29])
         );
  DFFARX1 \regf_reg[2][28]  ( .D(n139), .CLK(clk), .RSTB(n2305), .Q(reg3[28])
         );
  DFFARX1 \regf_reg[2][27]  ( .D(n138), .CLK(clk), .RSTB(n2304), .Q(reg3[27])
         );
  DFFARX1 \regf_reg[2][26]  ( .D(n137), .CLK(clk), .RSTB(n2304), .Q(reg3[26])
         );
  DFFARX1 \regf_reg[2][25]  ( .D(n136), .CLK(clk), .RSTB(n2304), .Q(reg3[25])
         );
  DFFARX1 \regf_reg[2][24]  ( .D(n135), .CLK(clk), .RSTB(n2304), .Q(reg3[24])
         );
  DFFARX1 \regf_reg[2][23]  ( .D(n134), .CLK(clk), .RSTB(n2304), .Q(reg3[23])
         );
  DFFARX1 \regf_reg[2][22]  ( .D(n133), .CLK(clk), .RSTB(n2304), .Q(reg3[22])
         );
  DFFARX1 \regf_reg[2][21]  ( .D(n132), .CLK(clk), .RSTB(n2304), .Q(reg3[21])
         );
  DFFARX1 \regf_reg[2][20]  ( .D(n131), .CLK(clk), .RSTB(n2304), .Q(reg3[20])
         );
  DFFARX1 \regf_reg[2][19]  ( .D(n130), .CLK(clk), .RSTB(n2304), .Q(reg3[19])
         );
  DFFARX1 \regf_reg[2][18]  ( .D(n129), .CLK(clk), .RSTB(n2304), .Q(reg3[18])
         );
  DFFARX1 \regf_reg[2][17]  ( .D(n128), .CLK(clk), .RSTB(n2304), .Q(reg3[17])
         );
  DFFARX1 \regf_reg[2][16]  ( .D(n127), .CLK(clk), .RSTB(n2304), .Q(reg3[16])
         );
  DFFARX1 \regf_reg[2][15]  ( .D(n126), .CLK(clk), .RSTB(n2303), .Q(reg3[15])
         );
  DFFARX1 \regf_reg[2][14]  ( .D(n125), .CLK(clk), .RSTB(n2303), .Q(reg3[14])
         );
  DFFARX1 \regf_reg[2][13]  ( .D(n124), .CLK(clk), .RSTB(n2303), .Q(reg3[13])
         );
  DFFARX1 \regf_reg[2][12]  ( .D(n123), .CLK(clk), .RSTB(n2303), .Q(reg3[12])
         );
  DFFARX1 \regf_reg[2][11]  ( .D(n122), .CLK(clk), .RSTB(n2303), .Q(reg3[11])
         );
  DFFARX1 \regf_reg[2][10]  ( .D(n121), .CLK(clk), .RSTB(n2303), .Q(reg3[10])
         );
  DFFARX1 \regf_reg[2][9]  ( .D(n120), .CLK(clk), .RSTB(n2303), .Q(reg3[9]) );
  DFFARX1 \regf_reg[2][8]  ( .D(n119), .CLK(clk), .RSTB(n2303), .Q(reg3[8]) );
  DFFARX1 \regf_reg[2][7]  ( .D(n118), .CLK(clk), .RSTB(n2303), .Q(reg3[7]) );
  DFFARX1 \regf_reg[2][6]  ( .D(n117), .CLK(clk), .RSTB(n2303), .Q(reg3[6]) );
  DFFARX1 \regf_reg[2][5]  ( .D(n116), .CLK(clk), .RSTB(n2303), .Q(reg3[5]) );
  DFFARX1 \regf_reg[2][4]  ( .D(n115), .CLK(clk), .RSTB(n2303), .Q(reg3[4]) );
  DFFARX1 \regf_reg[2][3]  ( .D(n114), .CLK(clk), .RSTB(n2302), .Q(reg3[3]) );
  DFFARX1 \regf_reg[2][2]  ( .D(n113), .CLK(clk), .RSTB(n2302), .Q(reg3[2]) );
  DFFARX1 \regf_reg[2][1]  ( .D(n112), .CLK(clk), .RSTB(n2302), .Q(reg3[1]) );
  DFFARX1 \regf_reg[2][0]  ( .D(n111), .CLK(clk), .RSTB(n2302), .Q(reg3[0]) );
  DFFARX1 \regf_reg[1][31]  ( .D(n110), .CLK(clk), .RSTB(n2302), .Q(reg2[31])
         );
  DFFARX1 \regf_reg[1][30]  ( .D(n109), .CLK(clk), .RSTB(n2302), .Q(reg2[30])
         );
  DFFARX1 \regf_reg[1][29]  ( .D(n108), .CLK(clk), .RSTB(n2302), .Q(reg2[29])
         );
  DFFARX1 \regf_reg[1][28]  ( .D(n107), .CLK(clk), .RSTB(n2302), .Q(reg2[28])
         );
  DFFARX1 \regf_reg[1][27]  ( .D(n106), .CLK(clk), .RSTB(n2302), .Q(reg2[27])
         );
  DFFARX1 \regf_reg[1][26]  ( .D(n105), .CLK(clk), .RSTB(n2302), .Q(reg2[26])
         );
  DFFARX1 \regf_reg[1][25]  ( .D(n104), .CLK(clk), .RSTB(n2302), .Q(reg2[25])
         );
  DFFARX1 \regf_reg[1][24]  ( .D(n103), .CLK(clk), .RSTB(n2302), .Q(reg2[24])
         );
  DFFARX1 \regf_reg[1][23]  ( .D(n102), .CLK(clk), .RSTB(n2301), .Q(reg2[23])
         );
  DFFARX1 \regf_reg[1][22]  ( .D(n101), .CLK(clk), .RSTB(n2301), .Q(reg2[22])
         );
  DFFARX1 \regf_reg[1][21]  ( .D(n100), .CLK(clk), .RSTB(n2301), .Q(reg2[21])
         );
  DFFARX1 \regf_reg[1][20]  ( .D(n99), .CLK(clk), .RSTB(n2301), .Q(reg2[20])
         );
  DFFARX1 \regf_reg[1][19]  ( .D(n98), .CLK(clk), .RSTB(n2301), .Q(reg2[19])
         );
  DFFARX1 \regf_reg[1][18]  ( .D(n97), .CLK(clk), .RSTB(n2301), .Q(reg2[18])
         );
  DFFARX1 \regf_reg[1][17]  ( .D(n96), .CLK(clk), .RSTB(n2301), .Q(reg2[17])
         );
  DFFARX1 \regf_reg[1][16]  ( .D(n95), .CLK(clk), .RSTB(n2301), .Q(reg2[16])
         );
  DFFARX1 \regf_reg[1][15]  ( .D(n94), .CLK(clk), .RSTB(n2301), .Q(reg2[15])
         );
  DFFARX1 \regf_reg[1][14]  ( .D(n93), .CLK(clk), .RSTB(n2301), .Q(reg2[14])
         );
  DFFARX1 \regf_reg[1][13]  ( .D(n92), .CLK(clk), .RSTB(n2301), .Q(reg2[13])
         );
  DFFARX1 \regf_reg[1][12]  ( .D(n91), .CLK(clk), .RSTB(n2301), .Q(reg2[12])
         );
  DFFARX1 \regf_reg[1][11]  ( .D(n90), .CLK(clk), .RSTB(n2300), .Q(reg2[11])
         );
  DFFARX1 \regf_reg[1][10]  ( .D(n89), .CLK(clk), .RSTB(n2300), .Q(reg2[10])
         );
  DFFARX1 \regf_reg[1][9]  ( .D(n88), .CLK(clk), .RSTB(n2300), .Q(reg2[9]) );
  DFFARX1 \regf_reg[1][8]  ( .D(n87), .CLK(clk), .RSTB(n2300), .Q(reg2[8]) );
  DFFARX1 \regf_reg[1][7]  ( .D(n86), .CLK(clk), .RSTB(n2300), .Q(reg2[7]) );
  DFFARX1 \regf_reg[1][6]  ( .D(n85), .CLK(clk), .RSTB(n2300), .Q(reg2[6]) );
  DFFARX1 \regf_reg[1][5]  ( .D(n84), .CLK(clk), .RSTB(n2300), .Q(reg2[5]) );
  DFFARX1 \regf_reg[1][4]  ( .D(n83), .CLK(clk), .RSTB(n2300), .Q(reg2[4]) );
  DFFARX1 \regf_reg[1][3]  ( .D(n82), .CLK(clk), .RSTB(n2300), .Q(reg2[3]) );
  DFFARX1 \regf_reg[1][2]  ( .D(n81), .CLK(clk), .RSTB(n2300), .Q(reg2[2]) );
  DFFARX1 \regf_reg[1][1]  ( .D(n80), .CLK(clk), .RSTB(n2300), .Q(reg2[1]) );
  DFFARX1 \regf_reg[1][0]  ( .D(n79), .CLK(clk), .RSTB(n2300), .Q(reg2[0]) );
  AO22X1 U100 ( .IN1(n2204), .IN2(n2203), .IN3(reg2[0]), .IN4(n37), .Q(n79) );
  AO22X1 U101 ( .IN1(n2207), .IN2(n2202), .IN3(reg2[1]), .IN4(n37), .Q(n80) );
  AO22X1 U102 ( .IN1(n2210), .IN2(n2203), .IN3(reg2[2]), .IN4(n37), .Q(n81) );
  AO22X1 U103 ( .IN1(n2213), .IN2(n2202), .IN3(reg2[3]), .IN4(n37), .Q(n82) );
  AO22X1 U104 ( .IN1(n2216), .IN2(n2202), .IN3(reg2[4]), .IN4(n37), .Q(n83) );
  AO22X1 U105 ( .IN1(n2219), .IN2(n2203), .IN3(reg2[5]), .IN4(n37), .Q(n84) );
  AO22X1 U106 ( .IN1(n2222), .IN2(n2202), .IN3(reg2[6]), .IN4(n37), .Q(n85) );
  AO22X1 U107 ( .IN1(n2225), .IN2(n2202), .IN3(reg2[7]), .IN4(n37), .Q(n86) );
  AO22X1 U108 ( .IN1(n2228), .IN2(n2203), .IN3(reg2[8]), .IN4(n2201), .Q(n87)
         );
  AO22X1 U109 ( .IN1(n2231), .IN2(n2203), .IN3(reg2[9]), .IN4(n2201), .Q(n88)
         );
  AO22X1 U110 ( .IN1(n2234), .IN2(n2202), .IN3(reg2[10]), .IN4(n2201), .Q(n89)
         );
  AO22X1 U111 ( .IN1(n2237), .IN2(n2202), .IN3(reg2[11]), .IN4(n2201), .Q(n90)
         );
  AO22X1 U112 ( .IN1(n2240), .IN2(n2202), .IN3(reg2[12]), .IN4(n2201), .Q(n91)
         );
  AO22X1 U113 ( .IN1(n2243), .IN2(n2202), .IN3(reg2[13]), .IN4(n2201), .Q(n92)
         );
  AO22X1 U114 ( .IN1(n2246), .IN2(n2202), .IN3(reg2[14]), .IN4(n2201), .Q(n93)
         );
  AO22X1 U115 ( .IN1(n2249), .IN2(n2202), .IN3(reg2[15]), .IN4(n2201), .Q(n94)
         );
  AO22X1 U116 ( .IN1(n2252), .IN2(n2202), .IN3(reg2[16]), .IN4(n2201), .Q(n95)
         );
  AO22X1 U117 ( .IN1(n2255), .IN2(n2202), .IN3(reg2[17]), .IN4(n2201), .Q(n96)
         );
  AO22X1 U118 ( .IN1(n2258), .IN2(n2203), .IN3(reg2[18]), .IN4(n2201), .Q(n97)
         );
  AO22X1 U119 ( .IN1(n2261), .IN2(n2202), .IN3(reg2[19]), .IN4(n2201), .Q(n98)
         );
  AO22X1 U120 ( .IN1(n2264), .IN2(n2203), .IN3(reg2[20]), .IN4(n2200), .Q(n99)
         );
  AO22X1 U121 ( .IN1(n2267), .IN2(n2202), .IN3(reg2[21]), .IN4(n2200), .Q(n100) );
  AO22X1 U122 ( .IN1(n2270), .IN2(n2203), .IN3(reg2[22]), .IN4(n2200), .Q(n101) );
  AO22X1 U123 ( .IN1(n2273), .IN2(n2202), .IN3(reg2[23]), .IN4(n2200), .Q(n102) );
  AO22X1 U124 ( .IN1(n2276), .IN2(n2203), .IN3(reg2[24]), .IN4(n2200), .Q(n103) );
  AO22X1 U125 ( .IN1(n2279), .IN2(n2203), .IN3(reg2[25]), .IN4(n2200), .Q(n104) );
  AO22X1 U126 ( .IN1(n2282), .IN2(n2203), .IN3(reg2[26]), .IN4(n2200), .Q(n105) );
  AO22X1 U127 ( .IN1(n2285), .IN2(n2203), .IN3(reg2[27]), .IN4(n2200), .Q(n106) );
  AO22X1 U128 ( .IN1(n2288), .IN2(n2203), .IN3(reg2[28]), .IN4(n2200), .Q(n107) );
  AO22X1 U129 ( .IN1(n2291), .IN2(n2203), .IN3(reg2[29]), .IN4(n2200), .Q(n108) );
  AO22X1 U130 ( .IN1(n2294), .IN2(n2203), .IN3(reg2[30]), .IN4(n2200), .Q(n109) );
  AO22X1 U131 ( .IN1(n2297), .IN2(n2203), .IN3(reg2[31]), .IN4(n2200), .Q(n110) );
  AO22X1 U132 ( .IN1(n2199), .IN2(n2204), .IN3(reg3[0]), .IN4(n40), .Q(n111)
         );
  AO22X1 U133 ( .IN1(n2198), .IN2(n2207), .IN3(reg3[1]), .IN4(n40), .Q(n112)
         );
  AO22X1 U134 ( .IN1(n2199), .IN2(n2210), .IN3(reg3[2]), .IN4(n40), .Q(n113)
         );
  AO22X1 U135 ( .IN1(n2198), .IN2(n2213), .IN3(reg3[3]), .IN4(n40), .Q(n114)
         );
  AO22X1 U136 ( .IN1(n2198), .IN2(n2216), .IN3(reg3[4]), .IN4(n40), .Q(n115)
         );
  AO22X1 U137 ( .IN1(n2199), .IN2(n2219), .IN3(reg3[5]), .IN4(n40), .Q(n116)
         );
  AO22X1 U138 ( .IN1(n2199), .IN2(n2222), .IN3(reg3[6]), .IN4(n40), .Q(n117)
         );
  AO22X1 U139 ( .IN1(n2198), .IN2(n2225), .IN3(reg3[7]), .IN4(n40), .Q(n118)
         );
  AO22X1 U140 ( .IN1(n2199), .IN2(n2228), .IN3(reg3[8]), .IN4(n2197), .Q(n119)
         );
  AO22X1 U141 ( .IN1(n2199), .IN2(n2231), .IN3(reg3[9]), .IN4(n2197), .Q(n120)
         );
  AO22X1 U142 ( .IN1(n2198), .IN2(n2234), .IN3(reg3[10]), .IN4(n2197), .Q(n121) );
  AO22X1 U143 ( .IN1(n2198), .IN2(n2237), .IN3(reg3[11]), .IN4(n2197), .Q(n122) );
  AO22X1 U144 ( .IN1(n2198), .IN2(n2240), .IN3(reg3[12]), .IN4(n2197), .Q(n123) );
  AO22X1 U145 ( .IN1(n2198), .IN2(n2243), .IN3(reg3[13]), .IN4(n2197), .Q(n124) );
  AO22X1 U146 ( .IN1(n2198), .IN2(n2246), .IN3(reg3[14]), .IN4(n2197), .Q(n125) );
  AO22X1 U147 ( .IN1(n2198), .IN2(n2249), .IN3(reg3[15]), .IN4(n2197), .Q(n126) );
  AO22X1 U148 ( .IN1(n2198), .IN2(n2252), .IN3(reg3[16]), .IN4(n2197), .Q(n127) );
  AO22X1 U149 ( .IN1(n2198), .IN2(n2255), .IN3(reg3[17]), .IN4(n2197), .Q(n128) );
  AO22X1 U150 ( .IN1(n2198), .IN2(n2258), .IN3(reg3[18]), .IN4(n2197), .Q(n129) );
  AO22X1 U151 ( .IN1(n2199), .IN2(n2261), .IN3(reg3[19]), .IN4(n2197), .Q(n130) );
  AO22X1 U152 ( .IN1(n2198), .IN2(n2264), .IN3(reg3[20]), .IN4(n2196), .Q(n131) );
  AO22X1 U153 ( .IN1(n2199), .IN2(n2267), .IN3(reg3[21]), .IN4(n2196), .Q(n132) );
  AO22X1 U154 ( .IN1(n2198), .IN2(n2270), .IN3(reg3[22]), .IN4(n2196), .Q(n133) );
  AO22X1 U155 ( .IN1(n2199), .IN2(n2273), .IN3(reg3[23]), .IN4(n2196), .Q(n134) );
  AO22X1 U156 ( .IN1(n2198), .IN2(n2276), .IN3(reg3[24]), .IN4(n2196), .Q(n135) );
  AO22X1 U157 ( .IN1(n2199), .IN2(n2279), .IN3(reg3[25]), .IN4(n2196), .Q(n136) );
  AO22X1 U158 ( .IN1(n2199), .IN2(n2282), .IN3(reg3[26]), .IN4(n2196), .Q(n137) );
  AO22X1 U159 ( .IN1(n2199), .IN2(n2285), .IN3(reg3[27]), .IN4(n2196), .Q(n138) );
  AO22X1 U160 ( .IN1(n2199), .IN2(n2288), .IN3(reg3[28]), .IN4(n2196), .Q(n139) );
  AO22X1 U161 ( .IN1(n2199), .IN2(n2291), .IN3(reg3[29]), .IN4(n2196), .Q(n140) );
  AO22X1 U162 ( .IN1(n2199), .IN2(n2294), .IN3(reg3[30]), .IN4(n2196), .Q(n141) );
  AO22X1 U163 ( .IN1(n2199), .IN2(n2297), .IN3(reg3[31]), .IN4(n2196), .Q(n142) );
  AO22X1 U164 ( .IN1(n2195), .IN2(n2204), .IN3(reg4[0]), .IN4(n42), .Q(n143)
         );
  AO22X1 U165 ( .IN1(n2194), .IN2(n2207), .IN3(reg4[1]), .IN4(n42), .Q(n144)
         );
  AO22X1 U166 ( .IN1(n2195), .IN2(n2210), .IN3(reg4[2]), .IN4(n42), .Q(n145)
         );
  AO22X1 U167 ( .IN1(n2194), .IN2(n2213), .IN3(reg4[3]), .IN4(n42), .Q(n146)
         );
  AO22X1 U168 ( .IN1(n2194), .IN2(n2216), .IN3(reg4[4]), .IN4(n42), .Q(n147)
         );
  AO22X1 U169 ( .IN1(n2195), .IN2(n2219), .IN3(reg4[5]), .IN4(n42), .Q(n148)
         );
  AO22X1 U170 ( .IN1(n2195), .IN2(n2222), .IN3(reg4[6]), .IN4(n42), .Q(n149)
         );
  AO22X1 U171 ( .IN1(n2194), .IN2(n2225), .IN3(reg4[7]), .IN4(n42), .Q(n150)
         );
  AO22X1 U172 ( .IN1(n2195), .IN2(n2228), .IN3(reg4[8]), .IN4(n2193), .Q(n151)
         );
  AO22X1 U173 ( .IN1(n2195), .IN2(n2231), .IN3(reg4[9]), .IN4(n2193), .Q(n152)
         );
  AO22X1 U174 ( .IN1(n2194), .IN2(n2234), .IN3(reg4[10]), .IN4(n2193), .Q(n153) );
  AO22X1 U175 ( .IN1(n2194), .IN2(n2237), .IN3(reg4[11]), .IN4(n2193), .Q(n154) );
  AO22X1 U176 ( .IN1(n2194), .IN2(n2240), .IN3(reg4[12]), .IN4(n2193), .Q(n155) );
  AO22X1 U177 ( .IN1(n2194), .IN2(n2243), .IN3(reg4[13]), .IN4(n2193), .Q(n156) );
  AO22X1 U178 ( .IN1(n2194), .IN2(n2246), .IN3(reg4[14]), .IN4(n2193), .Q(n157) );
  AO22X1 U179 ( .IN1(n2194), .IN2(n2249), .IN3(reg4[15]), .IN4(n2193), .Q(n158) );
  AO22X1 U180 ( .IN1(n2194), .IN2(n2252), .IN3(reg4[16]), .IN4(n2193), .Q(n159) );
  AO22X1 U181 ( .IN1(n2194), .IN2(n2255), .IN3(reg4[17]), .IN4(n2193), .Q(n160) );
  AO22X1 U182 ( .IN1(n2194), .IN2(n2258), .IN3(reg4[18]), .IN4(n2193), .Q(n161) );
  AO22X1 U183 ( .IN1(n2195), .IN2(n2261), .IN3(reg4[19]), .IN4(n2193), .Q(n162) );
  AO22X1 U184 ( .IN1(n2194), .IN2(n2264), .IN3(reg4[20]), .IN4(n2192), .Q(n163) );
  AO22X1 U185 ( .IN1(n2195), .IN2(n2267), .IN3(reg4[21]), .IN4(n2192), .Q(n164) );
  AO22X1 U186 ( .IN1(n2194), .IN2(n2270), .IN3(reg4[22]), .IN4(n2192), .Q(n165) );
  AO22X1 U187 ( .IN1(n2195), .IN2(n2273), .IN3(reg4[23]), .IN4(n2192), .Q(n166) );
  AO22X1 U188 ( .IN1(n2194), .IN2(n2276), .IN3(reg4[24]), .IN4(n2192), .Q(n167) );
  AO22X1 U189 ( .IN1(n2195), .IN2(n2279), .IN3(reg4[25]), .IN4(n2192), .Q(n168) );
  AO22X1 U190 ( .IN1(n2195), .IN2(n2282), .IN3(reg4[26]), .IN4(n2192), .Q(n169) );
  AO22X1 U191 ( .IN1(n2195), .IN2(n2285), .IN3(reg4[27]), .IN4(n2192), .Q(n170) );
  AO22X1 U192 ( .IN1(n2195), .IN2(n2288), .IN3(reg4[28]), .IN4(n2192), .Q(n171) );
  AO22X1 U193 ( .IN1(n2195), .IN2(n2291), .IN3(reg4[29]), .IN4(n2192), .Q(n172) );
  AO22X1 U194 ( .IN1(n2195), .IN2(n2294), .IN3(reg4[30]), .IN4(n2192), .Q(n173) );
  AO22X1 U195 ( .IN1(n2195), .IN2(n2297), .IN3(reg4[31]), .IN4(n2192), .Q(n174) );
  AO22X1 U196 ( .IN1(n2191), .IN2(n2204), .IN3(reg5[0]), .IN4(n44), .Q(n175)
         );
  AO22X1 U197 ( .IN1(n2190), .IN2(n2207), .IN3(reg5[1]), .IN4(n44), .Q(n176)
         );
  AO22X1 U198 ( .IN1(n2191), .IN2(n2210), .IN3(reg5[2]), .IN4(n44), .Q(n177)
         );
  AO22X1 U199 ( .IN1(n2190), .IN2(n2213), .IN3(reg5[3]), .IN4(n44), .Q(n178)
         );
  AO22X1 U200 ( .IN1(n2190), .IN2(n2216), .IN3(reg5[4]), .IN4(n44), .Q(n179)
         );
  AO22X1 U201 ( .IN1(n2191), .IN2(n2219), .IN3(reg5[5]), .IN4(n44), .Q(n180)
         );
  AO22X1 U202 ( .IN1(n2191), .IN2(n2222), .IN3(reg5[6]), .IN4(n44), .Q(n181)
         );
  AO22X1 U203 ( .IN1(n2190), .IN2(n2225), .IN3(reg5[7]), .IN4(n44), .Q(n182)
         );
  AO22X1 U204 ( .IN1(n2191), .IN2(n2228), .IN3(reg5[8]), .IN4(n2189), .Q(n183)
         );
  AO22X1 U205 ( .IN1(n2191), .IN2(n2231), .IN3(reg5[9]), .IN4(n2189), .Q(n184)
         );
  AO22X1 U206 ( .IN1(n2190), .IN2(n2234), .IN3(reg5[10]), .IN4(n2189), .Q(n185) );
  AO22X1 U207 ( .IN1(n2190), .IN2(n2237), .IN3(reg5[11]), .IN4(n2189), .Q(n186) );
  AO22X1 U208 ( .IN1(n2190), .IN2(n2240), .IN3(reg5[12]), .IN4(n2189), .Q(n187) );
  AO22X1 U209 ( .IN1(n2190), .IN2(n2243), .IN3(reg5[13]), .IN4(n2189), .Q(n188) );
  AO22X1 U210 ( .IN1(n2190), .IN2(n2246), .IN3(reg5[14]), .IN4(n2189), .Q(n189) );
  AO22X1 U211 ( .IN1(n2190), .IN2(n2249), .IN3(reg5[15]), .IN4(n2189), .Q(n190) );
  AO22X1 U212 ( .IN1(n2190), .IN2(n2252), .IN3(reg5[16]), .IN4(n2189), .Q(n191) );
  AO22X1 U213 ( .IN1(n2190), .IN2(n2255), .IN3(reg5[17]), .IN4(n2189), .Q(n192) );
  AO22X1 U214 ( .IN1(n2190), .IN2(n2258), .IN3(reg5[18]), .IN4(n2189), .Q(n193) );
  AO22X1 U215 ( .IN1(n2191), .IN2(n2261), .IN3(reg5[19]), .IN4(n2189), .Q(n194) );
  AO22X1 U216 ( .IN1(n2190), .IN2(n2264), .IN3(reg5[20]), .IN4(n2188), .Q(n195) );
  AO22X1 U217 ( .IN1(n2191), .IN2(n2267), .IN3(reg5[21]), .IN4(n2188), .Q(n196) );
  AO22X1 U218 ( .IN1(n2190), .IN2(n2270), .IN3(reg5[22]), .IN4(n2188), .Q(n197) );
  AO22X1 U219 ( .IN1(n2191), .IN2(n2273), .IN3(reg5[23]), .IN4(n2188), .Q(n198) );
  AO22X1 U220 ( .IN1(n2190), .IN2(n2276), .IN3(reg5[24]), .IN4(n2188), .Q(n199) );
  AO22X1 U221 ( .IN1(n2191), .IN2(n2279), .IN3(reg5[25]), .IN4(n2188), .Q(n200) );
  AO22X1 U222 ( .IN1(n2191), .IN2(n2282), .IN3(reg5[26]), .IN4(n2188), .Q(n201) );
  AO22X1 U223 ( .IN1(n2191), .IN2(n2285), .IN3(reg5[27]), .IN4(n2188), .Q(n202) );
  AO22X1 U224 ( .IN1(n2191), .IN2(n2288), .IN3(reg5[28]), .IN4(n2188), .Q(n203) );
  AO22X1 U225 ( .IN1(n2191), .IN2(n2291), .IN3(reg5[29]), .IN4(n2188), .Q(n204) );
  AO22X1 U226 ( .IN1(n2191), .IN2(n2294), .IN3(reg5[30]), .IN4(n2188), .Q(n205) );
  AO22X1 U227 ( .IN1(n2191), .IN2(n2297), .IN3(reg5[31]), .IN4(n2188), .Q(n206) );
  AO22X1 U228 ( .IN1(n2187), .IN2(n2204), .IN3(reg6[0]), .IN4(n46), .Q(n207)
         );
  AO22X1 U229 ( .IN1(n2186), .IN2(n2207), .IN3(reg6[1]), .IN4(n46), .Q(n208)
         );
  AO22X1 U230 ( .IN1(n2187), .IN2(n2210), .IN3(reg6[2]), .IN4(n46), .Q(n209)
         );
  AO22X1 U231 ( .IN1(n2186), .IN2(n2213), .IN3(reg6[3]), .IN4(n46), .Q(n210)
         );
  AO22X1 U232 ( .IN1(n2186), .IN2(n2216), .IN3(reg6[4]), .IN4(n46), .Q(n211)
         );
  AO22X1 U233 ( .IN1(n2187), .IN2(n2219), .IN3(reg6[5]), .IN4(n46), .Q(n212)
         );
  AO22X1 U234 ( .IN1(n2187), .IN2(n2222), .IN3(reg6[6]), .IN4(n46), .Q(n213)
         );
  AO22X1 U235 ( .IN1(n2186), .IN2(n2225), .IN3(reg6[7]), .IN4(n46), .Q(n214)
         );
  AO22X1 U236 ( .IN1(n2187), .IN2(n2228), .IN3(reg6[8]), .IN4(n2185), .Q(n215)
         );
  AO22X1 U237 ( .IN1(n2187), .IN2(n2231), .IN3(reg6[9]), .IN4(n2185), .Q(n216)
         );
  AO22X1 U238 ( .IN1(n2186), .IN2(n2234), .IN3(reg6[10]), .IN4(n2185), .Q(n217) );
  AO22X1 U239 ( .IN1(n2186), .IN2(n2237), .IN3(reg6[11]), .IN4(n2185), .Q(n218) );
  AO22X1 U240 ( .IN1(n2186), .IN2(n2240), .IN3(reg6[12]), .IN4(n2185), .Q(n219) );
  AO22X1 U241 ( .IN1(n2186), .IN2(n2243), .IN3(reg6[13]), .IN4(n2185), .Q(n220) );
  AO22X1 U242 ( .IN1(n2186), .IN2(n2246), .IN3(reg6[14]), .IN4(n2185), .Q(n221) );
  AO22X1 U243 ( .IN1(n2186), .IN2(n2249), .IN3(reg6[15]), .IN4(n2185), .Q(n222) );
  AO22X1 U244 ( .IN1(n2186), .IN2(n2252), .IN3(reg6[16]), .IN4(n2185), .Q(n223) );
  AO22X1 U245 ( .IN1(n2186), .IN2(n2255), .IN3(reg6[17]), .IN4(n2185), .Q(n224) );
  AO22X1 U246 ( .IN1(n2186), .IN2(n2258), .IN3(reg6[18]), .IN4(n2185), .Q(n225) );
  AO22X1 U247 ( .IN1(n2187), .IN2(n2261), .IN3(reg6[19]), .IN4(n2185), .Q(n226) );
  AO22X1 U248 ( .IN1(n2186), .IN2(n2264), .IN3(reg6[20]), .IN4(n2184), .Q(n227) );
  AO22X1 U249 ( .IN1(n2187), .IN2(n2267), .IN3(reg6[21]), .IN4(n2184), .Q(n228) );
  AO22X1 U250 ( .IN1(n2186), .IN2(n2270), .IN3(reg6[22]), .IN4(n2184), .Q(n229) );
  AO22X1 U251 ( .IN1(n2187), .IN2(n2273), .IN3(reg6[23]), .IN4(n2184), .Q(n230) );
  AO22X1 U252 ( .IN1(n2186), .IN2(n2276), .IN3(reg6[24]), .IN4(n2184), .Q(n231) );
  AO22X1 U253 ( .IN1(n2187), .IN2(n2279), .IN3(reg6[25]), .IN4(n2184), .Q(n232) );
  AO22X1 U254 ( .IN1(n2187), .IN2(n2282), .IN3(reg6[26]), .IN4(n2184), .Q(n233) );
  AO22X1 U255 ( .IN1(n2187), .IN2(n2285), .IN3(reg6[27]), .IN4(n2184), .Q(n234) );
  AO22X1 U256 ( .IN1(n2187), .IN2(n2288), .IN3(reg6[28]), .IN4(n2184), .Q(n235) );
  AO22X1 U257 ( .IN1(n2187), .IN2(n2291), .IN3(reg6[29]), .IN4(n2184), .Q(n236) );
  AO22X1 U258 ( .IN1(n2187), .IN2(n2294), .IN3(reg6[30]), .IN4(n2184), .Q(n237) );
  AO22X1 U259 ( .IN1(n2187), .IN2(n2297), .IN3(reg6[31]), .IN4(n2184), .Q(n238) );
  AO22X1 U260 ( .IN1(n2183), .IN2(n2204), .IN3(reg7[0]), .IN4(n48), .Q(n239)
         );
  AO22X1 U261 ( .IN1(n2182), .IN2(n2207), .IN3(reg7[1]), .IN4(n48), .Q(n240)
         );
  AO22X1 U262 ( .IN1(n2183), .IN2(n2210), .IN3(reg7[2]), .IN4(n48), .Q(n241)
         );
  AO22X1 U263 ( .IN1(n2182), .IN2(n2213), .IN3(reg7[3]), .IN4(n48), .Q(n242)
         );
  AO22X1 U264 ( .IN1(n2182), .IN2(n2216), .IN3(reg7[4]), .IN4(n48), .Q(n243)
         );
  AO22X1 U265 ( .IN1(n2183), .IN2(n2219), .IN3(reg7[5]), .IN4(n48), .Q(n244)
         );
  AO22X1 U266 ( .IN1(n2183), .IN2(n2222), .IN3(reg7[6]), .IN4(n48), .Q(n245)
         );
  AO22X1 U267 ( .IN1(n2182), .IN2(n2225), .IN3(reg7[7]), .IN4(n48), .Q(n246)
         );
  AO22X1 U268 ( .IN1(n2183), .IN2(n2228), .IN3(reg7[8]), .IN4(n2181), .Q(n247)
         );
  AO22X1 U269 ( .IN1(n2183), .IN2(n2231), .IN3(reg7[9]), .IN4(n2181), .Q(n248)
         );
  AO22X1 U270 ( .IN1(n2182), .IN2(n2234), .IN3(reg7[10]), .IN4(n2181), .Q(n249) );
  AO22X1 U271 ( .IN1(n2182), .IN2(n2237), .IN3(reg7[11]), .IN4(n2181), .Q(n250) );
  AO22X1 U272 ( .IN1(n2182), .IN2(n2240), .IN3(reg7[12]), .IN4(n2181), .Q(n251) );
  AO22X1 U273 ( .IN1(n2182), .IN2(n2243), .IN3(reg7[13]), .IN4(n2181), .Q(n252) );
  AO22X1 U274 ( .IN1(n2182), .IN2(n2246), .IN3(reg7[14]), .IN4(n2181), .Q(n253) );
  AO22X1 U275 ( .IN1(n2182), .IN2(n2249), .IN3(reg7[15]), .IN4(n2181), .Q(n254) );
  AO22X1 U276 ( .IN1(n2182), .IN2(n2252), .IN3(reg7[16]), .IN4(n2181), .Q(n255) );
  AO22X1 U277 ( .IN1(n2182), .IN2(n2255), .IN3(reg7[17]), .IN4(n2181), .Q(n256) );
  AO22X1 U278 ( .IN1(n2182), .IN2(n2258), .IN3(reg7[18]), .IN4(n2181), .Q(n257) );
  AO22X1 U279 ( .IN1(n2183), .IN2(n2261), .IN3(reg7[19]), .IN4(n2181), .Q(n258) );
  AO22X1 U280 ( .IN1(n2182), .IN2(n2264), .IN3(reg7[20]), .IN4(n2180), .Q(n259) );
  AO22X1 U281 ( .IN1(n2183), .IN2(n2267), .IN3(reg7[21]), .IN4(n2180), .Q(n260) );
  AO22X1 U282 ( .IN1(n2182), .IN2(n2270), .IN3(reg7[22]), .IN4(n2180), .Q(n261) );
  AO22X1 U283 ( .IN1(n2183), .IN2(n2273), .IN3(reg7[23]), .IN4(n2180), .Q(n262) );
  AO22X1 U284 ( .IN1(n2182), .IN2(n2276), .IN3(reg7[24]), .IN4(n2180), .Q(n263) );
  AO22X1 U285 ( .IN1(n2183), .IN2(n2279), .IN3(reg7[25]), .IN4(n2180), .Q(n264) );
  AO22X1 U286 ( .IN1(n2183), .IN2(n2282), .IN3(reg7[26]), .IN4(n2180), .Q(n265) );
  AO22X1 U287 ( .IN1(n2183), .IN2(n2285), .IN3(reg7[27]), .IN4(n2180), .Q(n266) );
  AO22X1 U288 ( .IN1(n2183), .IN2(n2288), .IN3(reg7[28]), .IN4(n2180), .Q(n267) );
  AO22X1 U289 ( .IN1(n2183), .IN2(n2291), .IN3(reg7[29]), .IN4(n2180), .Q(n268) );
  AO22X1 U290 ( .IN1(n2183), .IN2(n2294), .IN3(reg7[30]), .IN4(n2180), .Q(n269) );
  AO22X1 U291 ( .IN1(n2183), .IN2(n2297), .IN3(reg7[31]), .IN4(n2180), .Q(n270) );
  AO22X1 U292 ( .IN1(n2179), .IN2(n2204), .IN3(reg8[0]), .IN4(n50), .Q(n271)
         );
  AO22X1 U293 ( .IN1(n2178), .IN2(n2207), .IN3(reg8[1]), .IN4(n50), .Q(n272)
         );
  AO22X1 U294 ( .IN1(n2179), .IN2(n2210), .IN3(reg8[2]), .IN4(n50), .Q(n273)
         );
  AO22X1 U295 ( .IN1(n2178), .IN2(n2213), .IN3(reg8[3]), .IN4(n50), .Q(n274)
         );
  AO22X1 U296 ( .IN1(n2178), .IN2(n2216), .IN3(reg8[4]), .IN4(n50), .Q(n275)
         );
  AO22X1 U297 ( .IN1(n2179), .IN2(n2219), .IN3(reg8[5]), .IN4(n50), .Q(n276)
         );
  AO22X1 U298 ( .IN1(n2179), .IN2(n2222), .IN3(reg8[6]), .IN4(n50), .Q(n277)
         );
  AO22X1 U299 ( .IN1(n2178), .IN2(n2225), .IN3(reg8[7]), .IN4(n50), .Q(n278)
         );
  AO22X1 U300 ( .IN1(n2179), .IN2(n2228), .IN3(reg8[8]), .IN4(n2177), .Q(n279)
         );
  AO22X1 U301 ( .IN1(n2179), .IN2(n2231), .IN3(reg8[9]), .IN4(n2177), .Q(n280)
         );
  AO22X1 U302 ( .IN1(n2178), .IN2(n2234), .IN3(reg8[10]), .IN4(n2177), .Q(n281) );
  AO22X1 U303 ( .IN1(n2178), .IN2(n2237), .IN3(reg8[11]), .IN4(n2177), .Q(n282) );
  AO22X1 U304 ( .IN1(n2178), .IN2(n2240), .IN3(reg8[12]), .IN4(n2177), .Q(n283) );
  AO22X1 U305 ( .IN1(n2178), .IN2(n2243), .IN3(reg8[13]), .IN4(n2177), .Q(n284) );
  AO22X1 U306 ( .IN1(n2178), .IN2(n2246), .IN3(reg8[14]), .IN4(n2177), .Q(n285) );
  AO22X1 U307 ( .IN1(n2178), .IN2(n2249), .IN3(reg8[15]), .IN4(n2177), .Q(n286) );
  AO22X1 U308 ( .IN1(n2178), .IN2(n2252), .IN3(reg8[16]), .IN4(n2177), .Q(n287) );
  AO22X1 U309 ( .IN1(n2178), .IN2(n2255), .IN3(reg8[17]), .IN4(n2177), .Q(n288) );
  AO22X1 U310 ( .IN1(n2178), .IN2(n2258), .IN3(reg8[18]), .IN4(n2177), .Q(n289) );
  AO22X1 U311 ( .IN1(n2179), .IN2(n2261), .IN3(reg8[19]), .IN4(n2177), .Q(n290) );
  AO22X1 U312 ( .IN1(n2178), .IN2(n2264), .IN3(reg8[20]), .IN4(n2176), .Q(n291) );
  AO22X1 U313 ( .IN1(n2179), .IN2(n2267), .IN3(reg8[21]), .IN4(n2176), .Q(n292) );
  AO22X1 U314 ( .IN1(n2178), .IN2(n2270), .IN3(reg8[22]), .IN4(n2176), .Q(n293) );
  AO22X1 U315 ( .IN1(n2179), .IN2(n2273), .IN3(reg8[23]), .IN4(n2176), .Q(n294) );
  AO22X1 U316 ( .IN1(n2178), .IN2(n2276), .IN3(reg8[24]), .IN4(n2176), .Q(n295) );
  AO22X1 U317 ( .IN1(n2179), .IN2(n2279), .IN3(reg8[25]), .IN4(n2176), .Q(n296) );
  AO22X1 U318 ( .IN1(n2179), .IN2(n2282), .IN3(reg8[26]), .IN4(n2176), .Q(n297) );
  AO22X1 U319 ( .IN1(n2179), .IN2(n2285), .IN3(reg8[27]), .IN4(n2176), .Q(n298) );
  AO22X1 U320 ( .IN1(n2179), .IN2(n2288), .IN3(reg8[28]), .IN4(n2176), .Q(n299) );
  AO22X1 U321 ( .IN1(n2179), .IN2(n2291), .IN3(reg8[29]), .IN4(n2176), .Q(n300) );
  AO22X1 U322 ( .IN1(n2179), .IN2(n2294), .IN3(reg8[30]), .IN4(n2176), .Q(n301) );
  AO22X1 U323 ( .IN1(n2179), .IN2(n2297), .IN3(reg8[31]), .IN4(n2176), .Q(n302) );
  AND3X1 U324 ( .IN1(n2392), .IN2(n2393), .IN3(wr_en), .Q(n39) );
  AO22X1 U325 ( .IN1(n2175), .IN2(n2204), .IN3(reg9[0]), .IN4(n52), .Q(n303)
         );
  AO22X1 U326 ( .IN1(n2174), .IN2(n2207), .IN3(reg9[1]), .IN4(n52), .Q(n304)
         );
  AO22X1 U327 ( .IN1(n2175), .IN2(n2210), .IN3(reg9[2]), .IN4(n52), .Q(n305)
         );
  AO22X1 U328 ( .IN1(n2174), .IN2(n2213), .IN3(reg9[3]), .IN4(n52), .Q(n306)
         );
  AO22X1 U329 ( .IN1(n2174), .IN2(n2216), .IN3(reg9[4]), .IN4(n52), .Q(n307)
         );
  AO22X1 U330 ( .IN1(n2175), .IN2(n2219), .IN3(reg9[5]), .IN4(n52), .Q(n308)
         );
  AO22X1 U331 ( .IN1(n2175), .IN2(n2222), .IN3(reg9[6]), .IN4(n52), .Q(n309)
         );
  AO22X1 U332 ( .IN1(n2174), .IN2(n2225), .IN3(reg9[7]), .IN4(n52), .Q(n310)
         );
  AO22X1 U333 ( .IN1(n2175), .IN2(n2228), .IN3(reg9[8]), .IN4(n2173), .Q(n311)
         );
  AO22X1 U334 ( .IN1(n2175), .IN2(n2231), .IN3(reg9[9]), .IN4(n2173), .Q(n312)
         );
  AO22X1 U335 ( .IN1(n2174), .IN2(n2234), .IN3(reg9[10]), .IN4(n2173), .Q(n313) );
  AO22X1 U336 ( .IN1(n2174), .IN2(n2237), .IN3(reg9[11]), .IN4(n2173), .Q(n314) );
  AO22X1 U337 ( .IN1(n2174), .IN2(n2240), .IN3(reg9[12]), .IN4(n2173), .Q(n315) );
  AO22X1 U338 ( .IN1(n2174), .IN2(n2243), .IN3(reg9[13]), .IN4(n2173), .Q(n316) );
  AO22X1 U339 ( .IN1(n2174), .IN2(n2246), .IN3(reg9[14]), .IN4(n2173), .Q(n317) );
  AO22X1 U340 ( .IN1(n2174), .IN2(n2249), .IN3(reg9[15]), .IN4(n2173), .Q(n318) );
  AO22X1 U341 ( .IN1(n2174), .IN2(n2252), .IN3(reg9[16]), .IN4(n2173), .Q(n319) );
  AO22X1 U342 ( .IN1(n2174), .IN2(n2255), .IN3(reg9[17]), .IN4(n2173), .Q(n320) );
  AO22X1 U343 ( .IN1(n2174), .IN2(n2258), .IN3(reg9[18]), .IN4(n2173), .Q(n321) );
  AO22X1 U344 ( .IN1(n2175), .IN2(n2261), .IN3(reg9[19]), .IN4(n2173), .Q(n322) );
  AO22X1 U345 ( .IN1(n2174), .IN2(n2264), .IN3(reg9[20]), .IN4(n2172), .Q(n323) );
  AO22X1 U346 ( .IN1(n2175), .IN2(n2267), .IN3(reg9[21]), .IN4(n2172), .Q(n324) );
  AO22X1 U347 ( .IN1(n2174), .IN2(n2270), .IN3(reg9[22]), .IN4(n2172), .Q(n325) );
  AO22X1 U348 ( .IN1(n2175), .IN2(n2273), .IN3(reg9[23]), .IN4(n2172), .Q(n326) );
  AO22X1 U349 ( .IN1(n2174), .IN2(n2276), .IN3(reg9[24]), .IN4(n2172), .Q(n327) );
  AO22X1 U350 ( .IN1(n2175), .IN2(n2279), .IN3(reg9[25]), .IN4(n2172), .Q(n328) );
  AO22X1 U351 ( .IN1(n2175), .IN2(n2282), .IN3(reg9[26]), .IN4(n2172), .Q(n329) );
  AO22X1 U352 ( .IN1(n2175), .IN2(n2285), .IN3(reg9[27]), .IN4(n2172), .Q(n330) );
  AO22X1 U353 ( .IN1(n2175), .IN2(n2288), .IN3(reg9[28]), .IN4(n2172), .Q(n331) );
  AO22X1 U354 ( .IN1(n2175), .IN2(n2291), .IN3(reg9[29]), .IN4(n2172), .Q(n332) );
  AO22X1 U355 ( .IN1(n2175), .IN2(n2294), .IN3(reg9[30]), .IN4(n2172), .Q(n333) );
  AO22X1 U356 ( .IN1(n2175), .IN2(n2297), .IN3(reg9[31]), .IN4(n2172), .Q(n334) );
  AO22X1 U357 ( .IN1(n2171), .IN2(n2204), .IN3(reg10[0]), .IN4(n54), .Q(n335)
         );
  AO22X1 U358 ( .IN1(n2170), .IN2(n2207), .IN3(reg10[1]), .IN4(n54), .Q(n336)
         );
  AO22X1 U359 ( .IN1(n2171), .IN2(n2210), .IN3(reg10[2]), .IN4(n54), .Q(n337)
         );
  AO22X1 U360 ( .IN1(n2170), .IN2(n2213), .IN3(reg10[3]), .IN4(n54), .Q(n338)
         );
  AO22X1 U361 ( .IN1(n2170), .IN2(n2216), .IN3(reg10[4]), .IN4(n54), .Q(n339)
         );
  AO22X1 U362 ( .IN1(n2171), .IN2(n2219), .IN3(reg10[5]), .IN4(n54), .Q(n340)
         );
  AO22X1 U363 ( .IN1(n2171), .IN2(n2222), .IN3(reg10[6]), .IN4(n54), .Q(n341)
         );
  AO22X1 U364 ( .IN1(n2170), .IN2(n2225), .IN3(reg10[7]), .IN4(n54), .Q(n342)
         );
  AO22X1 U365 ( .IN1(n2171), .IN2(n2228), .IN3(reg10[8]), .IN4(n2169), .Q(n343) );
  AO22X1 U366 ( .IN1(n2171), .IN2(n2231), .IN3(reg10[9]), .IN4(n2169), .Q(n344) );
  AO22X1 U367 ( .IN1(n2170), .IN2(n2234), .IN3(reg10[10]), .IN4(n2169), .Q(
        n345) );
  AO22X1 U368 ( .IN1(n2170), .IN2(n2237), .IN3(reg10[11]), .IN4(n2169), .Q(
        n346) );
  AO22X1 U369 ( .IN1(n2170), .IN2(n2240), .IN3(reg10[12]), .IN4(n2169), .Q(
        n347) );
  AO22X1 U370 ( .IN1(n2170), .IN2(n2243), .IN3(reg10[13]), .IN4(n2169), .Q(
        n348) );
  AO22X1 U371 ( .IN1(n2170), .IN2(n2246), .IN3(reg10[14]), .IN4(n2169), .Q(
        n349) );
  AO22X1 U372 ( .IN1(n2170), .IN2(n2249), .IN3(reg10[15]), .IN4(n2169), .Q(
        n350) );
  AO22X1 U373 ( .IN1(n2170), .IN2(n2252), .IN3(reg10[16]), .IN4(n2169), .Q(
        n351) );
  AO22X1 U374 ( .IN1(n2170), .IN2(n2255), .IN3(reg10[17]), .IN4(n2169), .Q(
        n352) );
  AO22X1 U375 ( .IN1(n2170), .IN2(n2258), .IN3(reg10[18]), .IN4(n2169), .Q(
        n353) );
  AO22X1 U376 ( .IN1(n2171), .IN2(n2261), .IN3(reg10[19]), .IN4(n2169), .Q(
        n354) );
  AO22X1 U377 ( .IN1(n2170), .IN2(n2264), .IN3(reg10[20]), .IN4(n2168), .Q(
        n355) );
  AO22X1 U378 ( .IN1(n2171), .IN2(n2267), .IN3(reg10[21]), .IN4(n2168), .Q(
        n356) );
  AO22X1 U379 ( .IN1(n2170), .IN2(n2270), .IN3(reg10[22]), .IN4(n2168), .Q(
        n357) );
  AO22X1 U380 ( .IN1(n2171), .IN2(n2273), .IN3(reg10[23]), .IN4(n2168), .Q(
        n358) );
  AO22X1 U381 ( .IN1(n2170), .IN2(n2276), .IN3(reg10[24]), .IN4(n2168), .Q(
        n359) );
  AO22X1 U382 ( .IN1(n2171), .IN2(n2279), .IN3(reg10[25]), .IN4(n2168), .Q(
        n360) );
  AO22X1 U383 ( .IN1(n2171), .IN2(n2282), .IN3(reg10[26]), .IN4(n2168), .Q(
        n361) );
  AO22X1 U384 ( .IN1(n2171), .IN2(n2285), .IN3(reg10[27]), .IN4(n2168), .Q(
        n362) );
  AO22X1 U385 ( .IN1(n2171), .IN2(n2288), .IN3(reg10[28]), .IN4(n2168), .Q(
        n363) );
  AO22X1 U386 ( .IN1(n2171), .IN2(n2291), .IN3(reg10[29]), .IN4(n2168), .Q(
        n364) );
  AO22X1 U387 ( .IN1(n2171), .IN2(n2294), .IN3(reg10[30]), .IN4(n2168), .Q(
        n365) );
  AO22X1 U388 ( .IN1(n2171), .IN2(n2297), .IN3(reg10[31]), .IN4(n2168), .Q(
        n366) );
  AO22X1 U389 ( .IN1(n2167), .IN2(n2204), .IN3(reg11[0]), .IN4(n55), .Q(n367)
         );
  AO22X1 U390 ( .IN1(n2166), .IN2(n2207), .IN3(reg11[1]), .IN4(n55), .Q(n368)
         );
  AO22X1 U391 ( .IN1(n2167), .IN2(n2210), .IN3(reg11[2]), .IN4(n55), .Q(n369)
         );
  AO22X1 U392 ( .IN1(n2166), .IN2(n2213), .IN3(reg11[3]), .IN4(n55), .Q(n370)
         );
  AO22X1 U393 ( .IN1(n2166), .IN2(n2216), .IN3(reg11[4]), .IN4(n55), .Q(n371)
         );
  AO22X1 U394 ( .IN1(n2167), .IN2(n2219), .IN3(reg11[5]), .IN4(n55), .Q(n372)
         );
  AO22X1 U395 ( .IN1(n2167), .IN2(n2222), .IN3(reg11[6]), .IN4(n55), .Q(n373)
         );
  AO22X1 U396 ( .IN1(n2166), .IN2(n2225), .IN3(reg11[7]), .IN4(n55), .Q(n374)
         );
  AO22X1 U397 ( .IN1(n2167), .IN2(n2228), .IN3(reg11[8]), .IN4(n2165), .Q(n375) );
  AO22X1 U398 ( .IN1(n2167), .IN2(n2231), .IN3(reg11[9]), .IN4(n2165), .Q(n376) );
  AO22X1 U399 ( .IN1(n2166), .IN2(n2234), .IN3(reg11[10]), .IN4(n2165), .Q(
        n377) );
  AO22X1 U400 ( .IN1(n2166), .IN2(n2237), .IN3(reg11[11]), .IN4(n2165), .Q(
        n378) );
  AO22X1 U401 ( .IN1(n2166), .IN2(n2240), .IN3(reg11[12]), .IN4(n2165), .Q(
        n379) );
  AO22X1 U402 ( .IN1(n2166), .IN2(n2243), .IN3(reg11[13]), .IN4(n2165), .Q(
        n380) );
  AO22X1 U403 ( .IN1(n2166), .IN2(n2246), .IN3(reg11[14]), .IN4(n2165), .Q(
        n381) );
  AO22X1 U404 ( .IN1(n2166), .IN2(n2249), .IN3(reg11[15]), .IN4(n2165), .Q(
        n382) );
  AO22X1 U405 ( .IN1(n2166), .IN2(n2252), .IN3(reg11[16]), .IN4(n2165), .Q(
        n383) );
  AO22X1 U406 ( .IN1(n2166), .IN2(n2255), .IN3(reg11[17]), .IN4(n2165), .Q(
        n384) );
  AO22X1 U407 ( .IN1(n2166), .IN2(n2258), .IN3(reg11[18]), .IN4(n2165), .Q(
        n385) );
  AO22X1 U408 ( .IN1(n2167), .IN2(n2261), .IN3(reg11[19]), .IN4(n2165), .Q(
        n386) );
  AO22X1 U409 ( .IN1(n2166), .IN2(n2264), .IN3(reg11[20]), .IN4(n2164), .Q(
        n387) );
  AO22X1 U410 ( .IN1(n2167), .IN2(n2267), .IN3(reg11[21]), .IN4(n2164), .Q(
        n388) );
  AO22X1 U411 ( .IN1(n2166), .IN2(n2270), .IN3(reg11[22]), .IN4(n2164), .Q(
        n389) );
  AO22X1 U412 ( .IN1(n2167), .IN2(n2273), .IN3(reg11[23]), .IN4(n2164), .Q(
        n390) );
  AO22X1 U413 ( .IN1(n2166), .IN2(n2276), .IN3(reg11[24]), .IN4(n2164), .Q(
        n391) );
  AO22X1 U414 ( .IN1(n2167), .IN2(n2279), .IN3(reg11[25]), .IN4(n2164), .Q(
        n392) );
  AO22X1 U415 ( .IN1(n2167), .IN2(n2282), .IN3(reg11[26]), .IN4(n2164), .Q(
        n393) );
  AO22X1 U416 ( .IN1(n2167), .IN2(n2285), .IN3(reg11[27]), .IN4(n2164), .Q(
        n394) );
  AO22X1 U417 ( .IN1(n2167), .IN2(n2288), .IN3(reg11[28]), .IN4(n2164), .Q(
        n395) );
  AO22X1 U418 ( .IN1(n2167), .IN2(n2291), .IN3(reg11[29]), .IN4(n2164), .Q(
        n396) );
  AO22X1 U419 ( .IN1(n2167), .IN2(n2294), .IN3(reg11[30]), .IN4(n2164), .Q(
        n397) );
  AO22X1 U420 ( .IN1(n2167), .IN2(n2297), .IN3(reg11[31]), .IN4(n2164), .Q(
        n398) );
  AO22X1 U421 ( .IN1(n2163), .IN2(n2204), .IN3(reg12[0]), .IN4(n56), .Q(n399)
         );
  AO22X1 U422 ( .IN1(n2162), .IN2(n2207), .IN3(reg12[1]), .IN4(n56), .Q(n400)
         );
  AO22X1 U423 ( .IN1(n2163), .IN2(n2210), .IN3(reg12[2]), .IN4(n56), .Q(n401)
         );
  AO22X1 U424 ( .IN1(n2162), .IN2(n2213), .IN3(reg12[3]), .IN4(n56), .Q(n402)
         );
  AO22X1 U425 ( .IN1(n2162), .IN2(n2216), .IN3(reg12[4]), .IN4(n56), .Q(n403)
         );
  AO22X1 U426 ( .IN1(n2163), .IN2(n2219), .IN3(reg12[5]), .IN4(n56), .Q(n404)
         );
  AO22X1 U427 ( .IN1(n2163), .IN2(n2222), .IN3(reg12[6]), .IN4(n56), .Q(n405)
         );
  AO22X1 U428 ( .IN1(n2162), .IN2(n2225), .IN3(reg12[7]), .IN4(n56), .Q(n406)
         );
  AO22X1 U429 ( .IN1(n2163), .IN2(n2228), .IN3(reg12[8]), .IN4(n2161), .Q(n407) );
  AO22X1 U430 ( .IN1(n2163), .IN2(n2231), .IN3(reg12[9]), .IN4(n2161), .Q(n408) );
  AO22X1 U431 ( .IN1(n2162), .IN2(n2234), .IN3(reg12[10]), .IN4(n2161), .Q(
        n409) );
  AO22X1 U432 ( .IN1(n2162), .IN2(n2237), .IN3(reg12[11]), .IN4(n2161), .Q(
        n410) );
  AO22X1 U433 ( .IN1(n2162), .IN2(n2240), .IN3(reg12[12]), .IN4(n2161), .Q(
        n411) );
  AO22X1 U434 ( .IN1(n2162), .IN2(n2243), .IN3(reg12[13]), .IN4(n2161), .Q(
        n412) );
  AO22X1 U435 ( .IN1(n2162), .IN2(n2246), .IN3(reg12[14]), .IN4(n2161), .Q(
        n413) );
  AO22X1 U436 ( .IN1(n2162), .IN2(n2249), .IN3(reg12[15]), .IN4(n2161), .Q(
        n414) );
  AO22X1 U437 ( .IN1(n2162), .IN2(n2252), .IN3(reg12[16]), .IN4(n2161), .Q(
        n415) );
  AO22X1 U438 ( .IN1(n2162), .IN2(n2255), .IN3(reg12[17]), .IN4(n2161), .Q(
        n416) );
  AO22X1 U439 ( .IN1(n2162), .IN2(n2258), .IN3(reg12[18]), .IN4(n2161), .Q(
        n417) );
  AO22X1 U440 ( .IN1(n2163), .IN2(n2261), .IN3(reg12[19]), .IN4(n2161), .Q(
        n418) );
  AO22X1 U441 ( .IN1(n2162), .IN2(n2264), .IN3(reg12[20]), .IN4(n2160), .Q(
        n419) );
  AO22X1 U442 ( .IN1(n2163), .IN2(n2267), .IN3(reg12[21]), .IN4(n2160), .Q(
        n420) );
  AO22X1 U443 ( .IN1(n2162), .IN2(n2270), .IN3(reg12[22]), .IN4(n2160), .Q(
        n421) );
  AO22X1 U444 ( .IN1(n2163), .IN2(n2273), .IN3(reg12[23]), .IN4(n2160), .Q(
        n422) );
  AO22X1 U445 ( .IN1(n2162), .IN2(n2276), .IN3(reg12[24]), .IN4(n2160), .Q(
        n423) );
  AO22X1 U446 ( .IN1(n2163), .IN2(n2279), .IN3(reg12[25]), .IN4(n2160), .Q(
        n424) );
  AO22X1 U447 ( .IN1(n2163), .IN2(n2282), .IN3(reg12[26]), .IN4(n2160), .Q(
        n425) );
  AO22X1 U448 ( .IN1(n2163), .IN2(n2285), .IN3(reg12[27]), .IN4(n2160), .Q(
        n426) );
  AO22X1 U449 ( .IN1(n2163), .IN2(n2288), .IN3(reg12[28]), .IN4(n2160), .Q(
        n427) );
  AO22X1 U450 ( .IN1(n2163), .IN2(n2291), .IN3(reg12[29]), .IN4(n2160), .Q(
        n428) );
  AO22X1 U451 ( .IN1(n2163), .IN2(n2294), .IN3(reg12[30]), .IN4(n2160), .Q(
        n429) );
  AO22X1 U452 ( .IN1(n2163), .IN2(n2297), .IN3(reg12[31]), .IN4(n2160), .Q(
        n430) );
  AO22X1 U453 ( .IN1(n2159), .IN2(n2204), .IN3(reg13[0]), .IN4(n57), .Q(n431)
         );
  AO22X1 U454 ( .IN1(n2158), .IN2(n2207), .IN3(reg13[1]), .IN4(n57), .Q(n432)
         );
  AO22X1 U455 ( .IN1(n2159), .IN2(n2210), .IN3(reg13[2]), .IN4(n57), .Q(n433)
         );
  AO22X1 U456 ( .IN1(n2158), .IN2(n2213), .IN3(reg13[3]), .IN4(n57), .Q(n434)
         );
  AO22X1 U457 ( .IN1(n2158), .IN2(n2216), .IN3(reg13[4]), .IN4(n57), .Q(n435)
         );
  AO22X1 U458 ( .IN1(n2159), .IN2(n2219), .IN3(reg13[5]), .IN4(n57), .Q(n436)
         );
  AO22X1 U459 ( .IN1(n2159), .IN2(n2222), .IN3(reg13[6]), .IN4(n57), .Q(n437)
         );
  AO22X1 U460 ( .IN1(n2158), .IN2(n2225), .IN3(reg13[7]), .IN4(n57), .Q(n438)
         );
  AO22X1 U461 ( .IN1(n2159), .IN2(n2228), .IN3(reg13[8]), .IN4(n2157), .Q(n439) );
  AO22X1 U462 ( .IN1(n2159), .IN2(n2231), .IN3(reg13[9]), .IN4(n2157), .Q(n440) );
  AO22X1 U463 ( .IN1(n2158), .IN2(n2234), .IN3(reg13[10]), .IN4(n2157), .Q(
        n441) );
  AO22X1 U464 ( .IN1(n2158), .IN2(n2237), .IN3(reg13[11]), .IN4(n2157), .Q(
        n442) );
  AO22X1 U465 ( .IN1(n2158), .IN2(n2240), .IN3(reg13[12]), .IN4(n2157), .Q(
        n443) );
  AO22X1 U466 ( .IN1(n2158), .IN2(n2243), .IN3(reg13[13]), .IN4(n2157), .Q(
        n444) );
  AO22X1 U467 ( .IN1(n2158), .IN2(n2246), .IN3(reg13[14]), .IN4(n2157), .Q(
        n445) );
  AO22X1 U468 ( .IN1(n2158), .IN2(n2249), .IN3(reg13[15]), .IN4(n2157), .Q(
        n446) );
  AO22X1 U469 ( .IN1(n2158), .IN2(n2252), .IN3(reg13[16]), .IN4(n2157), .Q(
        n447) );
  AO22X1 U470 ( .IN1(n2158), .IN2(n2255), .IN3(reg13[17]), .IN4(n2157), .Q(
        n448) );
  AO22X1 U471 ( .IN1(n2158), .IN2(n2258), .IN3(reg13[18]), .IN4(n2157), .Q(
        n449) );
  AO22X1 U472 ( .IN1(n2159), .IN2(n2261), .IN3(reg13[19]), .IN4(n2157), .Q(
        n450) );
  AO22X1 U473 ( .IN1(n2158), .IN2(n2264), .IN3(reg13[20]), .IN4(n2156), .Q(
        n451) );
  AO22X1 U474 ( .IN1(n2159), .IN2(n2267), .IN3(reg13[21]), .IN4(n2156), .Q(
        n452) );
  AO22X1 U475 ( .IN1(n2158), .IN2(n2270), .IN3(reg13[22]), .IN4(n2156), .Q(
        n453) );
  AO22X1 U476 ( .IN1(n2159), .IN2(n2273), .IN3(reg13[23]), .IN4(n2156), .Q(
        n454) );
  AO22X1 U477 ( .IN1(n2158), .IN2(n2276), .IN3(reg13[24]), .IN4(n2156), .Q(
        n455) );
  AO22X1 U478 ( .IN1(n2159), .IN2(n2279), .IN3(reg13[25]), .IN4(n2156), .Q(
        n456) );
  AO22X1 U479 ( .IN1(n2159), .IN2(n2282), .IN3(reg13[26]), .IN4(n2156), .Q(
        n457) );
  AO22X1 U480 ( .IN1(n2159), .IN2(n2285), .IN3(reg13[27]), .IN4(n2156), .Q(
        n458) );
  AO22X1 U481 ( .IN1(n2159), .IN2(n2288), .IN3(reg13[28]), .IN4(n2156), .Q(
        n459) );
  AO22X1 U482 ( .IN1(n2159), .IN2(n2291), .IN3(reg13[29]), .IN4(n2156), .Q(
        n460) );
  AO22X1 U483 ( .IN1(n2159), .IN2(n2294), .IN3(reg13[30]), .IN4(n2156), .Q(
        n461) );
  AO22X1 U484 ( .IN1(n2159), .IN2(n2297), .IN3(reg13[31]), .IN4(n2156), .Q(
        n462) );
  AO22X1 U485 ( .IN1(n2155), .IN2(n2205), .IN3(reg14[0]), .IN4(n58), .Q(n463)
         );
  AO22X1 U486 ( .IN1(n2154), .IN2(n2208), .IN3(reg14[1]), .IN4(n58), .Q(n464)
         );
  AO22X1 U487 ( .IN1(n2155), .IN2(n2211), .IN3(reg14[2]), .IN4(n58), .Q(n465)
         );
  AO22X1 U488 ( .IN1(n2154), .IN2(n2214), .IN3(reg14[3]), .IN4(n58), .Q(n466)
         );
  AO22X1 U489 ( .IN1(n2154), .IN2(n2217), .IN3(reg14[4]), .IN4(n58), .Q(n467)
         );
  AO22X1 U490 ( .IN1(n2155), .IN2(n2220), .IN3(reg14[5]), .IN4(n58), .Q(n468)
         );
  AO22X1 U491 ( .IN1(n2155), .IN2(n2223), .IN3(reg14[6]), .IN4(n58), .Q(n469)
         );
  AO22X1 U492 ( .IN1(n2154), .IN2(n2226), .IN3(reg14[7]), .IN4(n58), .Q(n470)
         );
  AO22X1 U493 ( .IN1(n2155), .IN2(n2229), .IN3(reg14[8]), .IN4(n2153), .Q(n471) );
  AO22X1 U494 ( .IN1(n2155), .IN2(n2232), .IN3(reg14[9]), .IN4(n2153), .Q(n472) );
  AO22X1 U495 ( .IN1(n2154), .IN2(n2235), .IN3(reg14[10]), .IN4(n2153), .Q(
        n473) );
  AO22X1 U496 ( .IN1(n2154), .IN2(n2238), .IN3(reg14[11]), .IN4(n2153), .Q(
        n474) );
  AO22X1 U497 ( .IN1(n2154), .IN2(n2241), .IN3(reg14[12]), .IN4(n2153), .Q(
        n475) );
  AO22X1 U498 ( .IN1(n2154), .IN2(n2244), .IN3(reg14[13]), .IN4(n2153), .Q(
        n476) );
  AO22X1 U499 ( .IN1(n2154), .IN2(n2247), .IN3(reg14[14]), .IN4(n2153), .Q(
        n477) );
  AO22X1 U500 ( .IN1(n2154), .IN2(n2250), .IN3(reg14[15]), .IN4(n2153), .Q(
        n478) );
  AO22X1 U501 ( .IN1(n2154), .IN2(n2253), .IN3(reg14[16]), .IN4(n2153), .Q(
        n479) );
  AO22X1 U502 ( .IN1(n2154), .IN2(n2256), .IN3(reg14[17]), .IN4(n2153), .Q(
        n480) );
  AO22X1 U503 ( .IN1(n2154), .IN2(n2259), .IN3(reg14[18]), .IN4(n2153), .Q(
        n481) );
  AO22X1 U504 ( .IN1(n2155), .IN2(n2262), .IN3(reg14[19]), .IN4(n2153), .Q(
        n482) );
  AO22X1 U505 ( .IN1(n2154), .IN2(n2265), .IN3(reg14[20]), .IN4(n2152), .Q(
        n483) );
  AO22X1 U506 ( .IN1(n2155), .IN2(n2268), .IN3(reg14[21]), .IN4(n2152), .Q(
        n484) );
  AO22X1 U507 ( .IN1(n2154), .IN2(n2271), .IN3(reg14[22]), .IN4(n2152), .Q(
        n485) );
  AO22X1 U508 ( .IN1(n2155), .IN2(n2274), .IN3(reg14[23]), .IN4(n2152), .Q(
        n486) );
  AO22X1 U509 ( .IN1(n2154), .IN2(n2277), .IN3(reg14[24]), .IN4(n2152), .Q(
        n487) );
  AO22X1 U510 ( .IN1(n2155), .IN2(n2280), .IN3(reg14[25]), .IN4(n2152), .Q(
        n488) );
  AO22X1 U511 ( .IN1(n2155), .IN2(n2283), .IN3(reg14[26]), .IN4(n2152), .Q(
        n489) );
  AO22X1 U512 ( .IN1(n2155), .IN2(n2286), .IN3(reg14[27]), .IN4(n2152), .Q(
        n490) );
  AO22X1 U513 ( .IN1(n2155), .IN2(n2289), .IN3(reg14[28]), .IN4(n2152), .Q(
        n491) );
  AO22X1 U514 ( .IN1(n2155), .IN2(n2292), .IN3(reg14[29]), .IN4(n2152), .Q(
        n492) );
  AO22X1 U515 ( .IN1(n2155), .IN2(n2295), .IN3(reg14[30]), .IN4(n2152), .Q(
        n493) );
  AO22X1 U516 ( .IN1(n2155), .IN2(n2298), .IN3(reg14[31]), .IN4(n2152), .Q(
        n494) );
  AO22X1 U517 ( .IN1(n2151), .IN2(n2205), .IN3(reg15[0]), .IN4(n59), .Q(n495)
         );
  AO22X1 U518 ( .IN1(n2150), .IN2(n2208), .IN3(reg15[1]), .IN4(n59), .Q(n496)
         );
  AO22X1 U519 ( .IN1(n2151), .IN2(n2211), .IN3(reg15[2]), .IN4(n59), .Q(n497)
         );
  AO22X1 U520 ( .IN1(n2150), .IN2(n2214), .IN3(reg15[3]), .IN4(n59), .Q(n498)
         );
  AO22X1 U521 ( .IN1(n2150), .IN2(n2217), .IN3(reg15[4]), .IN4(n59), .Q(n499)
         );
  AO22X1 U522 ( .IN1(n2151), .IN2(n2220), .IN3(reg15[5]), .IN4(n59), .Q(n500)
         );
  AO22X1 U523 ( .IN1(n2151), .IN2(n2223), .IN3(reg15[6]), .IN4(n59), .Q(n501)
         );
  AO22X1 U524 ( .IN1(n2150), .IN2(n2226), .IN3(reg15[7]), .IN4(n59), .Q(n502)
         );
  AO22X1 U525 ( .IN1(n2151), .IN2(n2229), .IN3(reg15[8]), .IN4(n2149), .Q(n503) );
  AO22X1 U526 ( .IN1(n2151), .IN2(n2232), .IN3(reg15[9]), .IN4(n2149), .Q(n504) );
  AO22X1 U527 ( .IN1(n2150), .IN2(n2235), .IN3(reg15[10]), .IN4(n2149), .Q(
        n505) );
  AO22X1 U528 ( .IN1(n2150), .IN2(n2238), .IN3(reg15[11]), .IN4(n2149), .Q(
        n506) );
  AO22X1 U529 ( .IN1(n2150), .IN2(n2241), .IN3(reg15[12]), .IN4(n2149), .Q(
        n507) );
  AO22X1 U530 ( .IN1(n2150), .IN2(n2244), .IN3(reg15[13]), .IN4(n2149), .Q(
        n508) );
  AO22X1 U531 ( .IN1(n2150), .IN2(n2247), .IN3(reg15[14]), .IN4(n2149), .Q(
        n509) );
  AO22X1 U532 ( .IN1(n2150), .IN2(n2250), .IN3(reg15[15]), .IN4(n2149), .Q(
        n510) );
  AO22X1 U533 ( .IN1(n2150), .IN2(n2253), .IN3(reg15[16]), .IN4(n2149), .Q(
        n511) );
  AO22X1 U534 ( .IN1(n2150), .IN2(n2256), .IN3(reg15[17]), .IN4(n2149), .Q(
        n512) );
  AO22X1 U535 ( .IN1(n2150), .IN2(n2259), .IN3(reg15[18]), .IN4(n2149), .Q(
        n513) );
  AO22X1 U536 ( .IN1(n2151), .IN2(n2262), .IN3(reg15[19]), .IN4(n2149), .Q(
        n514) );
  AO22X1 U537 ( .IN1(n2150), .IN2(n2265), .IN3(reg15[20]), .IN4(n2148), .Q(
        n515) );
  AO22X1 U538 ( .IN1(n2151), .IN2(n2268), .IN3(reg15[21]), .IN4(n2148), .Q(
        n516) );
  AO22X1 U539 ( .IN1(n2150), .IN2(n2271), .IN3(reg15[22]), .IN4(n2148), .Q(
        n517) );
  AO22X1 U540 ( .IN1(n2151), .IN2(n2274), .IN3(reg15[23]), .IN4(n2148), .Q(
        n518) );
  AO22X1 U541 ( .IN1(n2150), .IN2(n2277), .IN3(reg15[24]), .IN4(n2148), .Q(
        n519) );
  AO22X1 U542 ( .IN1(n2151), .IN2(n2280), .IN3(reg15[25]), .IN4(n2148), .Q(
        n520) );
  AO22X1 U543 ( .IN1(n2151), .IN2(n2283), .IN3(reg15[26]), .IN4(n2148), .Q(
        n521) );
  AO22X1 U544 ( .IN1(n2151), .IN2(n2286), .IN3(reg15[27]), .IN4(n2148), .Q(
        n522) );
  AO22X1 U545 ( .IN1(n2151), .IN2(n2289), .IN3(reg15[28]), .IN4(n2148), .Q(
        n523) );
  AO22X1 U546 ( .IN1(n2151), .IN2(n2292), .IN3(reg15[29]), .IN4(n2148), .Q(
        n524) );
  AO22X1 U547 ( .IN1(n2151), .IN2(n2295), .IN3(reg15[30]), .IN4(n2148), .Q(
        n525) );
  AO22X1 U548 ( .IN1(n2151), .IN2(n2298), .IN3(reg15[31]), .IN4(n2148), .Q(
        n526) );
  AO22X1 U549 ( .IN1(n2147), .IN2(n2205), .IN3(reg16[0]), .IN4(n60), .Q(n527)
         );
  AO22X1 U550 ( .IN1(n2146), .IN2(n2208), .IN3(reg16[1]), .IN4(n60), .Q(n528)
         );
  AO22X1 U551 ( .IN1(n2147), .IN2(n2211), .IN3(reg16[2]), .IN4(n60), .Q(n529)
         );
  AO22X1 U552 ( .IN1(n2146), .IN2(n2214), .IN3(reg16[3]), .IN4(n60), .Q(n530)
         );
  AO22X1 U553 ( .IN1(n2146), .IN2(n2217), .IN3(reg16[4]), .IN4(n60), .Q(n531)
         );
  AO22X1 U554 ( .IN1(n2147), .IN2(n2220), .IN3(reg16[5]), .IN4(n60), .Q(n532)
         );
  AO22X1 U555 ( .IN1(n2147), .IN2(n2223), .IN3(reg16[6]), .IN4(n60), .Q(n533)
         );
  AO22X1 U556 ( .IN1(n2146), .IN2(n2226), .IN3(reg16[7]), .IN4(n60), .Q(n534)
         );
  AO22X1 U557 ( .IN1(n2147), .IN2(n2229), .IN3(reg16[8]), .IN4(n2145), .Q(n535) );
  AO22X1 U558 ( .IN1(n2147), .IN2(n2232), .IN3(reg16[9]), .IN4(n2145), .Q(n536) );
  AO22X1 U559 ( .IN1(n2146), .IN2(n2235), .IN3(reg16[10]), .IN4(n2145), .Q(
        n537) );
  AO22X1 U560 ( .IN1(n2146), .IN2(n2238), .IN3(reg16[11]), .IN4(n2145), .Q(
        n538) );
  AO22X1 U561 ( .IN1(n2146), .IN2(n2241), .IN3(reg16[12]), .IN4(n2145), .Q(
        n539) );
  AO22X1 U562 ( .IN1(n2146), .IN2(n2244), .IN3(reg16[13]), .IN4(n2145), .Q(
        n540) );
  AO22X1 U563 ( .IN1(n2146), .IN2(n2247), .IN3(reg16[14]), .IN4(n2145), .Q(
        n541) );
  AO22X1 U564 ( .IN1(n2146), .IN2(n2250), .IN3(reg16[15]), .IN4(n2145), .Q(
        n542) );
  AO22X1 U565 ( .IN1(n2146), .IN2(n2253), .IN3(reg16[16]), .IN4(n2145), .Q(
        n543) );
  AO22X1 U566 ( .IN1(n2146), .IN2(n2256), .IN3(reg16[17]), .IN4(n2145), .Q(
        n544) );
  AO22X1 U567 ( .IN1(n2146), .IN2(n2259), .IN3(reg16[18]), .IN4(n2145), .Q(
        n545) );
  AO22X1 U568 ( .IN1(n2147), .IN2(n2262), .IN3(reg16[19]), .IN4(n2145), .Q(
        n546) );
  AO22X1 U569 ( .IN1(n2146), .IN2(n2265), .IN3(reg16[20]), .IN4(n2144), .Q(
        n547) );
  AO22X1 U570 ( .IN1(n2147), .IN2(n2268), .IN3(reg16[21]), .IN4(n2144), .Q(
        n548) );
  AO22X1 U571 ( .IN1(n2146), .IN2(n2271), .IN3(reg16[22]), .IN4(n2144), .Q(
        n549) );
  AO22X1 U572 ( .IN1(n2147), .IN2(n2274), .IN3(reg16[23]), .IN4(n2144), .Q(
        n550) );
  AO22X1 U573 ( .IN1(n2146), .IN2(n2277), .IN3(reg16[24]), .IN4(n2144), .Q(
        n551) );
  AO22X1 U574 ( .IN1(n2147), .IN2(n2280), .IN3(reg16[25]), .IN4(n2144), .Q(
        n552) );
  AO22X1 U575 ( .IN1(n2147), .IN2(n2283), .IN3(reg16[26]), .IN4(n2144), .Q(
        n553) );
  AO22X1 U576 ( .IN1(n2147), .IN2(n2286), .IN3(reg16[27]), .IN4(n2144), .Q(
        n554) );
  AO22X1 U577 ( .IN1(n2147), .IN2(n2289), .IN3(reg16[28]), .IN4(n2144), .Q(
        n555) );
  AO22X1 U578 ( .IN1(n2147), .IN2(n2292), .IN3(reg16[29]), .IN4(n2144), .Q(
        n556) );
  AO22X1 U579 ( .IN1(n2147), .IN2(n2295), .IN3(reg16[30]), .IN4(n2144), .Q(
        n557) );
  AO22X1 U580 ( .IN1(n2147), .IN2(n2298), .IN3(reg16[31]), .IN4(n2144), .Q(
        n558) );
  AND3X1 U581 ( .IN1(wr_en), .IN2(n2393), .IN3(wr_addr[3]), .Q(n53) );
  AO22X1 U582 ( .IN1(n2143), .IN2(n2205), .IN3(reg17[0]), .IN4(n61), .Q(n559)
         );
  AO22X1 U583 ( .IN1(n2142), .IN2(n2208), .IN3(reg17[1]), .IN4(n61), .Q(n560)
         );
  AO22X1 U584 ( .IN1(n2143), .IN2(n2211), .IN3(reg17[2]), .IN4(n61), .Q(n561)
         );
  AO22X1 U585 ( .IN1(n2142), .IN2(n2214), .IN3(reg17[3]), .IN4(n61), .Q(n562)
         );
  AO22X1 U586 ( .IN1(n2142), .IN2(n2217), .IN3(reg17[4]), .IN4(n61), .Q(n563)
         );
  AO22X1 U587 ( .IN1(n2143), .IN2(n2220), .IN3(reg17[5]), .IN4(n61), .Q(n564)
         );
  AO22X1 U588 ( .IN1(n2143), .IN2(n2223), .IN3(reg17[6]), .IN4(n61), .Q(n565)
         );
  AO22X1 U589 ( .IN1(n2142), .IN2(n2226), .IN3(reg17[7]), .IN4(n61), .Q(n566)
         );
  AO22X1 U590 ( .IN1(n2143), .IN2(n2229), .IN3(reg17[8]), .IN4(n2141), .Q(n567) );
  AO22X1 U591 ( .IN1(n2143), .IN2(n2232), .IN3(reg17[9]), .IN4(n2141), .Q(n568) );
  AO22X1 U592 ( .IN1(n2142), .IN2(n2235), .IN3(reg17[10]), .IN4(n2141), .Q(
        n569) );
  AO22X1 U593 ( .IN1(n2142), .IN2(n2238), .IN3(reg17[11]), .IN4(n2141), .Q(
        n570) );
  AO22X1 U594 ( .IN1(n2142), .IN2(n2241), .IN3(reg17[12]), .IN4(n2141), .Q(
        n571) );
  AO22X1 U595 ( .IN1(n2142), .IN2(n2244), .IN3(reg17[13]), .IN4(n2141), .Q(
        n572) );
  AO22X1 U596 ( .IN1(n2142), .IN2(n2247), .IN3(reg17[14]), .IN4(n2141), .Q(
        n573) );
  AO22X1 U597 ( .IN1(n2142), .IN2(n2250), .IN3(reg17[15]), .IN4(n2141), .Q(
        n574) );
  AO22X1 U598 ( .IN1(n2142), .IN2(n2253), .IN3(reg17[16]), .IN4(n2141), .Q(
        n575) );
  AO22X1 U599 ( .IN1(n2142), .IN2(n2256), .IN3(reg17[17]), .IN4(n2141), .Q(
        n576) );
  AO22X1 U600 ( .IN1(n2142), .IN2(n2259), .IN3(reg17[18]), .IN4(n2141), .Q(
        n577) );
  AO22X1 U601 ( .IN1(n2143), .IN2(n2262), .IN3(reg17[19]), .IN4(n2141), .Q(
        n578) );
  AO22X1 U602 ( .IN1(n2142), .IN2(n2265), .IN3(reg17[20]), .IN4(n2140), .Q(
        n579) );
  AO22X1 U603 ( .IN1(n2143), .IN2(n2268), .IN3(reg17[21]), .IN4(n2140), .Q(
        n580) );
  AO22X1 U604 ( .IN1(n2142), .IN2(n2271), .IN3(reg17[22]), .IN4(n2140), .Q(
        n581) );
  AO22X1 U605 ( .IN1(n2143), .IN2(n2274), .IN3(reg17[23]), .IN4(n2140), .Q(
        n582) );
  AO22X1 U606 ( .IN1(n2142), .IN2(n2277), .IN3(reg17[24]), .IN4(n2140), .Q(
        n583) );
  AO22X1 U607 ( .IN1(n2143), .IN2(n2280), .IN3(reg17[25]), .IN4(n2140), .Q(
        n584) );
  AO22X1 U608 ( .IN1(n2143), .IN2(n2283), .IN3(reg17[26]), .IN4(n2140), .Q(
        n585) );
  AO22X1 U609 ( .IN1(n2143), .IN2(n2286), .IN3(reg17[27]), .IN4(n2140), .Q(
        n586) );
  AO22X1 U610 ( .IN1(n2143), .IN2(n2289), .IN3(reg17[28]), .IN4(n2140), .Q(
        n587) );
  AO22X1 U611 ( .IN1(n2143), .IN2(n2292), .IN3(reg17[29]), .IN4(n2140), .Q(
        n588) );
  AO22X1 U612 ( .IN1(n2143), .IN2(n2295), .IN3(reg17[30]), .IN4(n2140), .Q(
        n589) );
  AO22X1 U613 ( .IN1(n2143), .IN2(n2298), .IN3(reg17[31]), .IN4(n2140), .Q(
        n590) );
  AO22X1 U614 ( .IN1(n2139), .IN2(n2205), .IN3(reg18[0]), .IN4(n63), .Q(n591)
         );
  AO22X1 U615 ( .IN1(n2138), .IN2(n2208), .IN3(reg18[1]), .IN4(n63), .Q(n592)
         );
  AO22X1 U616 ( .IN1(n2139), .IN2(n2211), .IN3(reg18[2]), .IN4(n63), .Q(n593)
         );
  AO22X1 U617 ( .IN1(n2138), .IN2(n2214), .IN3(reg18[3]), .IN4(n63), .Q(n594)
         );
  AO22X1 U618 ( .IN1(n2138), .IN2(n2217), .IN3(reg18[4]), .IN4(n63), .Q(n595)
         );
  AO22X1 U619 ( .IN1(n2139), .IN2(n2220), .IN3(reg18[5]), .IN4(n63), .Q(n596)
         );
  AO22X1 U620 ( .IN1(n2139), .IN2(n2223), .IN3(reg18[6]), .IN4(n63), .Q(n597)
         );
  AO22X1 U621 ( .IN1(n2138), .IN2(n2226), .IN3(reg18[7]), .IN4(n63), .Q(n598)
         );
  AO22X1 U622 ( .IN1(n2139), .IN2(n2229), .IN3(reg18[8]), .IN4(n2137), .Q(n599) );
  AO22X1 U623 ( .IN1(n2139), .IN2(n2232), .IN3(reg18[9]), .IN4(n2137), .Q(n600) );
  AO22X1 U624 ( .IN1(n2138), .IN2(n2235), .IN3(reg18[10]), .IN4(n2137), .Q(
        n601) );
  AO22X1 U625 ( .IN1(n2138), .IN2(n2238), .IN3(reg18[11]), .IN4(n2137), .Q(
        n602) );
  AO22X1 U626 ( .IN1(n2138), .IN2(n2241), .IN3(reg18[12]), .IN4(n2137), .Q(
        n603) );
  AO22X1 U627 ( .IN1(n2138), .IN2(n2244), .IN3(reg18[13]), .IN4(n2137), .Q(
        n604) );
  AO22X1 U628 ( .IN1(n2138), .IN2(n2247), .IN3(reg18[14]), .IN4(n2137), .Q(
        n605) );
  AO22X1 U629 ( .IN1(n2138), .IN2(n2250), .IN3(reg18[15]), .IN4(n2137), .Q(
        n606) );
  AO22X1 U630 ( .IN1(n2138), .IN2(n2253), .IN3(reg18[16]), .IN4(n2137), .Q(
        n607) );
  AO22X1 U631 ( .IN1(n2138), .IN2(n2256), .IN3(reg18[17]), .IN4(n2137), .Q(
        n608) );
  AO22X1 U632 ( .IN1(n2138), .IN2(n2259), .IN3(reg18[18]), .IN4(n2137), .Q(
        n609) );
  AO22X1 U633 ( .IN1(n2139), .IN2(n2262), .IN3(reg18[19]), .IN4(n2137), .Q(
        n610) );
  AO22X1 U634 ( .IN1(n2138), .IN2(n2265), .IN3(reg18[20]), .IN4(n2136), .Q(
        n611) );
  AO22X1 U635 ( .IN1(n2139), .IN2(n2268), .IN3(reg18[21]), .IN4(n2136), .Q(
        n612) );
  AO22X1 U636 ( .IN1(n2138), .IN2(n2271), .IN3(reg18[22]), .IN4(n2136), .Q(
        n613) );
  AO22X1 U637 ( .IN1(n2139), .IN2(n2274), .IN3(reg18[23]), .IN4(n2136), .Q(
        n614) );
  AO22X1 U638 ( .IN1(n2138), .IN2(n2277), .IN3(reg18[24]), .IN4(n2136), .Q(
        n615) );
  AO22X1 U639 ( .IN1(n2139), .IN2(n2280), .IN3(reg18[25]), .IN4(n2136), .Q(
        n616) );
  AO22X1 U640 ( .IN1(n2139), .IN2(n2283), .IN3(reg18[26]), .IN4(n2136), .Q(
        n617) );
  AO22X1 U641 ( .IN1(n2139), .IN2(n2286), .IN3(reg18[27]), .IN4(n2136), .Q(
        n618) );
  AO22X1 U642 ( .IN1(n2139), .IN2(n2289), .IN3(reg18[28]), .IN4(n2136), .Q(
        n619) );
  AO22X1 U643 ( .IN1(n2139), .IN2(n2292), .IN3(reg18[29]), .IN4(n2136), .Q(
        n620) );
  AO22X1 U644 ( .IN1(n2139), .IN2(n2295), .IN3(reg18[30]), .IN4(n2136), .Q(
        n621) );
  AO22X1 U645 ( .IN1(n2139), .IN2(n2298), .IN3(reg18[31]), .IN4(n2136), .Q(
        n622) );
  AO22X1 U646 ( .IN1(n2135), .IN2(n2205), .IN3(reg19[0]), .IN4(n64), .Q(n623)
         );
  AO22X1 U647 ( .IN1(n2134), .IN2(n2208), .IN3(reg19[1]), .IN4(n64), .Q(n624)
         );
  AO22X1 U648 ( .IN1(n2135), .IN2(n2211), .IN3(reg19[2]), .IN4(n64), .Q(n625)
         );
  AO22X1 U649 ( .IN1(n2134), .IN2(n2214), .IN3(reg19[3]), .IN4(n64), .Q(n626)
         );
  AO22X1 U650 ( .IN1(n2134), .IN2(n2217), .IN3(reg19[4]), .IN4(n64), .Q(n627)
         );
  AO22X1 U651 ( .IN1(n2135), .IN2(n2220), .IN3(reg19[5]), .IN4(n64), .Q(n628)
         );
  AO22X1 U652 ( .IN1(n2135), .IN2(n2223), .IN3(reg19[6]), .IN4(n64), .Q(n629)
         );
  AO22X1 U653 ( .IN1(n2134), .IN2(n2226), .IN3(reg19[7]), .IN4(n64), .Q(n630)
         );
  AO22X1 U654 ( .IN1(n2135), .IN2(n2229), .IN3(reg19[8]), .IN4(n2133), .Q(n631) );
  AO22X1 U655 ( .IN1(n2135), .IN2(n2232), .IN3(reg19[9]), .IN4(n2133), .Q(n632) );
  AO22X1 U656 ( .IN1(n2134), .IN2(n2235), .IN3(reg19[10]), .IN4(n2133), .Q(
        n633) );
  AO22X1 U657 ( .IN1(n2134), .IN2(n2238), .IN3(reg19[11]), .IN4(n2133), .Q(
        n634) );
  AO22X1 U658 ( .IN1(n2134), .IN2(n2241), .IN3(reg19[12]), .IN4(n2133), .Q(
        n635) );
  AO22X1 U659 ( .IN1(n2134), .IN2(n2244), .IN3(reg19[13]), .IN4(n2133), .Q(
        n636) );
  AO22X1 U660 ( .IN1(n2134), .IN2(n2247), .IN3(reg19[14]), .IN4(n2133), .Q(
        n637) );
  AO22X1 U661 ( .IN1(n2134), .IN2(n2250), .IN3(reg19[15]), .IN4(n2133), .Q(
        n638) );
  AO22X1 U662 ( .IN1(n2134), .IN2(n2253), .IN3(reg19[16]), .IN4(n2133), .Q(
        n639) );
  AO22X1 U663 ( .IN1(n2134), .IN2(n2256), .IN3(reg19[17]), .IN4(n2133), .Q(
        n640) );
  AO22X1 U664 ( .IN1(n2134), .IN2(n2259), .IN3(reg19[18]), .IN4(n2133), .Q(
        n641) );
  AO22X1 U665 ( .IN1(n2135), .IN2(n2262), .IN3(reg19[19]), .IN4(n2133), .Q(
        n642) );
  AO22X1 U666 ( .IN1(n2134), .IN2(n2265), .IN3(reg19[20]), .IN4(n2132), .Q(
        n643) );
  AO22X1 U667 ( .IN1(n2135), .IN2(n2268), .IN3(reg19[21]), .IN4(n2132), .Q(
        n644) );
  AO22X1 U668 ( .IN1(n2134), .IN2(n2271), .IN3(reg19[22]), .IN4(n2132), .Q(
        n645) );
  AO22X1 U669 ( .IN1(n2135), .IN2(n2274), .IN3(reg19[23]), .IN4(n2132), .Q(
        n646) );
  AO22X1 U670 ( .IN1(n2134), .IN2(n2277), .IN3(reg19[24]), .IN4(n2132), .Q(
        n647) );
  AO22X1 U671 ( .IN1(n2135), .IN2(n2280), .IN3(reg19[25]), .IN4(n2132), .Q(
        n648) );
  AO22X1 U672 ( .IN1(n2135), .IN2(n2283), .IN3(reg19[26]), .IN4(n2132), .Q(
        n649) );
  AO22X1 U673 ( .IN1(n2135), .IN2(n2286), .IN3(reg19[27]), .IN4(n2132), .Q(
        n650) );
  AO22X1 U674 ( .IN1(n2135), .IN2(n2289), .IN3(reg19[28]), .IN4(n2132), .Q(
        n651) );
  AO22X1 U675 ( .IN1(n2135), .IN2(n2292), .IN3(reg19[29]), .IN4(n2132), .Q(
        n652) );
  AO22X1 U676 ( .IN1(n2135), .IN2(n2295), .IN3(reg19[30]), .IN4(n2132), .Q(
        n653) );
  AO22X1 U677 ( .IN1(n2135), .IN2(n2298), .IN3(reg19[31]), .IN4(n2132), .Q(
        n654) );
  AO22X1 U678 ( .IN1(n2131), .IN2(n2205), .IN3(reg20[0]), .IN4(n65), .Q(n655)
         );
  AO22X1 U679 ( .IN1(n2130), .IN2(n2208), .IN3(reg20[1]), .IN4(n65), .Q(n656)
         );
  AO22X1 U680 ( .IN1(n2131), .IN2(n2211), .IN3(reg20[2]), .IN4(n65), .Q(n657)
         );
  AO22X1 U681 ( .IN1(n2130), .IN2(n2214), .IN3(reg20[3]), .IN4(n65), .Q(n658)
         );
  AO22X1 U682 ( .IN1(n2130), .IN2(n2217), .IN3(reg20[4]), .IN4(n65), .Q(n659)
         );
  AO22X1 U683 ( .IN1(n2131), .IN2(n2220), .IN3(reg20[5]), .IN4(n65), .Q(n660)
         );
  AO22X1 U684 ( .IN1(n2131), .IN2(n2223), .IN3(reg20[6]), .IN4(n65), .Q(n661)
         );
  AO22X1 U685 ( .IN1(n2130), .IN2(n2226), .IN3(reg20[7]), .IN4(n65), .Q(n662)
         );
  AO22X1 U686 ( .IN1(n2131), .IN2(n2229), .IN3(reg20[8]), .IN4(n2129), .Q(n663) );
  AO22X1 U687 ( .IN1(n2131), .IN2(n2232), .IN3(reg20[9]), .IN4(n2129), .Q(n664) );
  AO22X1 U688 ( .IN1(n2130), .IN2(n2235), .IN3(reg20[10]), .IN4(n2129), .Q(
        n665) );
  AO22X1 U689 ( .IN1(n2130), .IN2(n2238), .IN3(reg20[11]), .IN4(n2129), .Q(
        n666) );
  AO22X1 U690 ( .IN1(n2130), .IN2(n2241), .IN3(reg20[12]), .IN4(n2129), .Q(
        n667) );
  AO22X1 U691 ( .IN1(n2130), .IN2(n2244), .IN3(reg20[13]), .IN4(n2129), .Q(
        n668) );
  AO22X1 U692 ( .IN1(n2130), .IN2(n2247), .IN3(reg20[14]), .IN4(n2129), .Q(
        n669) );
  AO22X1 U693 ( .IN1(n2130), .IN2(n2250), .IN3(reg20[15]), .IN4(n2129), .Q(
        n670) );
  AO22X1 U694 ( .IN1(n2130), .IN2(n2253), .IN3(reg20[16]), .IN4(n2129), .Q(
        n671) );
  AO22X1 U695 ( .IN1(n2130), .IN2(n2256), .IN3(reg20[17]), .IN4(n2129), .Q(
        n672) );
  AO22X1 U696 ( .IN1(n2130), .IN2(n2259), .IN3(reg20[18]), .IN4(n2129), .Q(
        n673) );
  AO22X1 U697 ( .IN1(n2131), .IN2(n2262), .IN3(reg20[19]), .IN4(n2129), .Q(
        n674) );
  AO22X1 U698 ( .IN1(n2130), .IN2(n2265), .IN3(reg20[20]), .IN4(n2128), .Q(
        n675) );
  AO22X1 U699 ( .IN1(n2131), .IN2(n2268), .IN3(reg20[21]), .IN4(n2128), .Q(
        n676) );
  AO22X1 U700 ( .IN1(n2130), .IN2(n2271), .IN3(reg20[22]), .IN4(n2128), .Q(
        n677) );
  AO22X1 U701 ( .IN1(n2131), .IN2(n2274), .IN3(reg20[23]), .IN4(n2128), .Q(
        n678) );
  AO22X1 U702 ( .IN1(n2130), .IN2(n2277), .IN3(reg20[24]), .IN4(n2128), .Q(
        n679) );
  AO22X1 U703 ( .IN1(n2131), .IN2(n2280), .IN3(reg20[25]), .IN4(n2128), .Q(
        n680) );
  AO22X1 U704 ( .IN1(n2131), .IN2(n2283), .IN3(reg20[26]), .IN4(n2128), .Q(
        n681) );
  AO22X1 U705 ( .IN1(n2131), .IN2(n2286), .IN3(reg20[27]), .IN4(n2128), .Q(
        n682) );
  AO22X1 U706 ( .IN1(n2131), .IN2(n2289), .IN3(reg20[28]), .IN4(n2128), .Q(
        n683) );
  AO22X1 U707 ( .IN1(n2131), .IN2(n2292), .IN3(reg20[29]), .IN4(n2128), .Q(
        n684) );
  AO22X1 U708 ( .IN1(n2131), .IN2(n2295), .IN3(reg20[30]), .IN4(n2128), .Q(
        n685) );
  AO22X1 U709 ( .IN1(n2131), .IN2(n2298), .IN3(reg20[31]), .IN4(n2128), .Q(
        n686) );
  AO22X1 U710 ( .IN1(n2127), .IN2(n2205), .IN3(reg21[0]), .IN4(n66), .Q(n687)
         );
  AO22X1 U711 ( .IN1(n2126), .IN2(n2208), .IN3(reg21[1]), .IN4(n66), .Q(n688)
         );
  AO22X1 U712 ( .IN1(n2127), .IN2(n2211), .IN3(reg21[2]), .IN4(n66), .Q(n689)
         );
  AO22X1 U713 ( .IN1(n2126), .IN2(n2214), .IN3(reg21[3]), .IN4(n66), .Q(n690)
         );
  AO22X1 U714 ( .IN1(n2126), .IN2(n2217), .IN3(reg21[4]), .IN4(n66), .Q(n691)
         );
  AO22X1 U715 ( .IN1(n2127), .IN2(n2220), .IN3(reg21[5]), .IN4(n66), .Q(n692)
         );
  AO22X1 U716 ( .IN1(n2127), .IN2(n2223), .IN3(reg21[6]), .IN4(n66), .Q(n693)
         );
  AO22X1 U717 ( .IN1(n2126), .IN2(n2226), .IN3(reg21[7]), .IN4(n66), .Q(n694)
         );
  AO22X1 U718 ( .IN1(n2127), .IN2(n2229), .IN3(reg21[8]), .IN4(n2125), .Q(n695) );
  AO22X1 U719 ( .IN1(n2127), .IN2(n2232), .IN3(reg21[9]), .IN4(n2125), .Q(n696) );
  AO22X1 U720 ( .IN1(n2126), .IN2(n2235), .IN3(reg21[10]), .IN4(n2125), .Q(
        n697) );
  AO22X1 U721 ( .IN1(n2126), .IN2(n2238), .IN3(reg21[11]), .IN4(n2125), .Q(
        n698) );
  AO22X1 U722 ( .IN1(n2126), .IN2(n2241), .IN3(reg21[12]), .IN4(n2125), .Q(
        n699) );
  AO22X1 U723 ( .IN1(n2126), .IN2(n2244), .IN3(reg21[13]), .IN4(n2125), .Q(
        n700) );
  AO22X1 U724 ( .IN1(n2126), .IN2(n2247), .IN3(reg21[14]), .IN4(n2125), .Q(
        n701) );
  AO22X1 U725 ( .IN1(n2126), .IN2(n2250), .IN3(reg21[15]), .IN4(n2125), .Q(
        n702) );
  AO22X1 U726 ( .IN1(n2126), .IN2(n2253), .IN3(reg21[16]), .IN4(n2125), .Q(
        n703) );
  AO22X1 U727 ( .IN1(n2126), .IN2(n2256), .IN3(reg21[17]), .IN4(n2125), .Q(
        n704) );
  AO22X1 U728 ( .IN1(n2126), .IN2(n2259), .IN3(reg21[18]), .IN4(n2125), .Q(
        n705) );
  AO22X1 U729 ( .IN1(n2127), .IN2(n2262), .IN3(reg21[19]), .IN4(n2125), .Q(
        n706) );
  AO22X1 U730 ( .IN1(n2126), .IN2(n2265), .IN3(reg21[20]), .IN4(n2124), .Q(
        n707) );
  AO22X1 U731 ( .IN1(n2127), .IN2(n2268), .IN3(reg21[21]), .IN4(n2124), .Q(
        n708) );
  AO22X1 U732 ( .IN1(n2126), .IN2(n2271), .IN3(reg21[22]), .IN4(n2124), .Q(
        n709) );
  AO22X1 U733 ( .IN1(n2127), .IN2(n2274), .IN3(reg21[23]), .IN4(n2124), .Q(
        n710) );
  AO22X1 U734 ( .IN1(n2126), .IN2(n2277), .IN3(reg21[24]), .IN4(n2124), .Q(
        n711) );
  AO22X1 U735 ( .IN1(n2127), .IN2(n2280), .IN3(reg21[25]), .IN4(n2124), .Q(
        n712) );
  AO22X1 U736 ( .IN1(n2127), .IN2(n2283), .IN3(reg21[26]), .IN4(n2124), .Q(
        n713) );
  AO22X1 U737 ( .IN1(n2127), .IN2(n2286), .IN3(reg21[27]), .IN4(n2124), .Q(
        n714) );
  AO22X1 U738 ( .IN1(n2127), .IN2(n2289), .IN3(reg21[28]), .IN4(n2124), .Q(
        n715) );
  AO22X1 U739 ( .IN1(n2127), .IN2(n2292), .IN3(reg21[29]), .IN4(n2124), .Q(
        n716) );
  AO22X1 U740 ( .IN1(n2127), .IN2(n2295), .IN3(reg21[30]), .IN4(n2124), .Q(
        n717) );
  AO22X1 U741 ( .IN1(n2127), .IN2(n2298), .IN3(reg21[31]), .IN4(n2124), .Q(
        n718) );
  AO22X1 U742 ( .IN1(n2123), .IN2(n2205), .IN3(reg22[0]), .IN4(n67), .Q(n719)
         );
  AO22X1 U743 ( .IN1(n2122), .IN2(n2208), .IN3(reg22[1]), .IN4(n67), .Q(n720)
         );
  AO22X1 U744 ( .IN1(n2123), .IN2(n2211), .IN3(reg22[2]), .IN4(n67), .Q(n721)
         );
  AO22X1 U745 ( .IN1(n2122), .IN2(n2214), .IN3(reg22[3]), .IN4(n67), .Q(n722)
         );
  AO22X1 U746 ( .IN1(n2122), .IN2(n2217), .IN3(reg22[4]), .IN4(n67), .Q(n723)
         );
  AO22X1 U747 ( .IN1(n2123), .IN2(n2220), .IN3(reg22[5]), .IN4(n67), .Q(n724)
         );
  AO22X1 U748 ( .IN1(n2123), .IN2(n2223), .IN3(reg22[6]), .IN4(n67), .Q(n725)
         );
  AO22X1 U749 ( .IN1(n2122), .IN2(n2226), .IN3(reg22[7]), .IN4(n67), .Q(n726)
         );
  AO22X1 U750 ( .IN1(n2123), .IN2(n2229), .IN3(reg22[8]), .IN4(n2121), .Q(n727) );
  AO22X1 U751 ( .IN1(n2123), .IN2(n2232), .IN3(reg22[9]), .IN4(n2121), .Q(n728) );
  AO22X1 U752 ( .IN1(n2122), .IN2(n2235), .IN3(reg22[10]), .IN4(n2121), .Q(
        n729) );
  AO22X1 U753 ( .IN1(n2122), .IN2(n2238), .IN3(reg22[11]), .IN4(n2121), .Q(
        n730) );
  AO22X1 U754 ( .IN1(n2122), .IN2(n2241), .IN3(reg22[12]), .IN4(n2121), .Q(
        n731) );
  AO22X1 U755 ( .IN1(n2122), .IN2(n2244), .IN3(reg22[13]), .IN4(n2121), .Q(
        n732) );
  AO22X1 U756 ( .IN1(n2122), .IN2(n2247), .IN3(reg22[14]), .IN4(n2121), .Q(
        n733) );
  AO22X1 U757 ( .IN1(n2122), .IN2(n2250), .IN3(reg22[15]), .IN4(n2121), .Q(
        n734) );
  AO22X1 U758 ( .IN1(n2122), .IN2(n2253), .IN3(reg22[16]), .IN4(n2121), .Q(
        n735) );
  AO22X1 U759 ( .IN1(n2122), .IN2(n2256), .IN3(reg22[17]), .IN4(n2121), .Q(
        n736) );
  AO22X1 U760 ( .IN1(n2122), .IN2(n2259), .IN3(reg22[18]), .IN4(n2121), .Q(
        n737) );
  AO22X1 U761 ( .IN1(n2123), .IN2(n2262), .IN3(reg22[19]), .IN4(n2121), .Q(
        n738) );
  AO22X1 U762 ( .IN1(n2122), .IN2(n2265), .IN3(reg22[20]), .IN4(n2120), .Q(
        n739) );
  AO22X1 U763 ( .IN1(n2123), .IN2(n2268), .IN3(reg22[21]), .IN4(n2120), .Q(
        n740) );
  AO22X1 U764 ( .IN1(n2122), .IN2(n2271), .IN3(reg22[22]), .IN4(n2120), .Q(
        n741) );
  AO22X1 U765 ( .IN1(n2123), .IN2(n2274), .IN3(reg22[23]), .IN4(n2120), .Q(
        n742) );
  AO22X1 U766 ( .IN1(n2122), .IN2(n2277), .IN3(reg22[24]), .IN4(n2120), .Q(
        n743) );
  AO22X1 U767 ( .IN1(n2123), .IN2(n2280), .IN3(reg22[25]), .IN4(n2120), .Q(
        n744) );
  AO22X1 U768 ( .IN1(n2123), .IN2(n2283), .IN3(reg22[26]), .IN4(n2120), .Q(
        n745) );
  AO22X1 U769 ( .IN1(n2123), .IN2(n2286), .IN3(reg22[27]), .IN4(n2120), .Q(
        n746) );
  AO22X1 U770 ( .IN1(n2123), .IN2(n2289), .IN3(reg22[28]), .IN4(n2120), .Q(
        n747) );
  AO22X1 U771 ( .IN1(n2123), .IN2(n2292), .IN3(reg22[29]), .IN4(n2120), .Q(
        n748) );
  AO22X1 U772 ( .IN1(n2123), .IN2(n2295), .IN3(reg22[30]), .IN4(n2120), .Q(
        n749) );
  AO22X1 U773 ( .IN1(n2123), .IN2(n2298), .IN3(reg22[31]), .IN4(n2120), .Q(
        n750) );
  AO22X1 U774 ( .IN1(n2119), .IN2(n2205), .IN3(reg23[0]), .IN4(n68), .Q(n751)
         );
  AO22X1 U775 ( .IN1(n2118), .IN2(n2208), .IN3(reg23[1]), .IN4(n68), .Q(n752)
         );
  AO22X1 U776 ( .IN1(n2119), .IN2(n2211), .IN3(reg23[2]), .IN4(n68), .Q(n753)
         );
  AO22X1 U777 ( .IN1(n2118), .IN2(n2214), .IN3(reg23[3]), .IN4(n68), .Q(n754)
         );
  AO22X1 U778 ( .IN1(n2118), .IN2(n2217), .IN3(reg23[4]), .IN4(n68), .Q(n755)
         );
  AO22X1 U779 ( .IN1(n2119), .IN2(n2220), .IN3(reg23[5]), .IN4(n68), .Q(n756)
         );
  AO22X1 U780 ( .IN1(n2119), .IN2(n2223), .IN3(reg23[6]), .IN4(n68), .Q(n757)
         );
  AO22X1 U781 ( .IN1(n2118), .IN2(n2226), .IN3(reg23[7]), .IN4(n68), .Q(n758)
         );
  AO22X1 U782 ( .IN1(n2119), .IN2(n2229), .IN3(reg23[8]), .IN4(n2117), .Q(n759) );
  AO22X1 U783 ( .IN1(n2119), .IN2(n2232), .IN3(reg23[9]), .IN4(n2117), .Q(n760) );
  AO22X1 U784 ( .IN1(n2118), .IN2(n2235), .IN3(reg23[10]), .IN4(n2117), .Q(
        n761) );
  AO22X1 U785 ( .IN1(n2118), .IN2(n2238), .IN3(reg23[11]), .IN4(n2117), .Q(
        n762) );
  AO22X1 U786 ( .IN1(n2118), .IN2(n2241), .IN3(reg23[12]), .IN4(n2117), .Q(
        n763) );
  AO22X1 U787 ( .IN1(n2118), .IN2(n2244), .IN3(reg23[13]), .IN4(n2117), .Q(
        n764) );
  AO22X1 U788 ( .IN1(n2118), .IN2(n2247), .IN3(reg23[14]), .IN4(n2117), .Q(
        n765) );
  AO22X1 U789 ( .IN1(n2118), .IN2(n2250), .IN3(reg23[15]), .IN4(n2117), .Q(
        n766) );
  AO22X1 U790 ( .IN1(n2118), .IN2(n2253), .IN3(reg23[16]), .IN4(n2117), .Q(
        n767) );
  AO22X1 U791 ( .IN1(n2118), .IN2(n2256), .IN3(reg23[17]), .IN4(n2117), .Q(
        n768) );
  AO22X1 U792 ( .IN1(n2118), .IN2(n2259), .IN3(reg23[18]), .IN4(n2117), .Q(
        n769) );
  AO22X1 U793 ( .IN1(n2119), .IN2(n2262), .IN3(reg23[19]), .IN4(n2117), .Q(
        n770) );
  AO22X1 U794 ( .IN1(n2118), .IN2(n2265), .IN3(reg23[20]), .IN4(n2116), .Q(
        n771) );
  AO22X1 U795 ( .IN1(n2119), .IN2(n2268), .IN3(reg23[21]), .IN4(n2116), .Q(
        n772) );
  AO22X1 U796 ( .IN1(n2118), .IN2(n2271), .IN3(reg23[22]), .IN4(n2116), .Q(
        n773) );
  AO22X1 U797 ( .IN1(n2119), .IN2(n2274), .IN3(reg23[23]), .IN4(n2116), .Q(
        n774) );
  AO22X1 U798 ( .IN1(n2118), .IN2(n2277), .IN3(reg23[24]), .IN4(n2116), .Q(
        n775) );
  AO22X1 U799 ( .IN1(n2119), .IN2(n2280), .IN3(reg23[25]), .IN4(n2116), .Q(
        n776) );
  AO22X1 U800 ( .IN1(n2119), .IN2(n2283), .IN3(reg23[26]), .IN4(n2116), .Q(
        n777) );
  AO22X1 U801 ( .IN1(n2119), .IN2(n2286), .IN3(reg23[27]), .IN4(n2116), .Q(
        n778) );
  AO22X1 U802 ( .IN1(n2119), .IN2(n2289), .IN3(reg23[28]), .IN4(n2116), .Q(
        n779) );
  AO22X1 U803 ( .IN1(n2119), .IN2(n2292), .IN3(reg23[29]), .IN4(n2116), .Q(
        n780) );
  AO22X1 U804 ( .IN1(n2119), .IN2(n2295), .IN3(reg23[30]), .IN4(n2116), .Q(
        n781) );
  AO22X1 U805 ( .IN1(n2119), .IN2(n2298), .IN3(reg23[31]), .IN4(n2116), .Q(
        n782) );
  AO22X1 U806 ( .IN1(n2115), .IN2(n2205), .IN3(reg24[0]), .IN4(n69), .Q(n783)
         );
  AO22X1 U807 ( .IN1(n2114), .IN2(n2208), .IN3(reg24[1]), .IN4(n69), .Q(n784)
         );
  AO22X1 U808 ( .IN1(n2115), .IN2(n2211), .IN3(reg24[2]), .IN4(n69), .Q(n785)
         );
  AO22X1 U809 ( .IN1(n2114), .IN2(n2214), .IN3(reg24[3]), .IN4(n69), .Q(n786)
         );
  AO22X1 U810 ( .IN1(n2114), .IN2(n2217), .IN3(reg24[4]), .IN4(n69), .Q(n787)
         );
  AO22X1 U811 ( .IN1(n2115), .IN2(n2220), .IN3(reg24[5]), .IN4(n69), .Q(n788)
         );
  AO22X1 U812 ( .IN1(n2115), .IN2(n2223), .IN3(reg24[6]), .IN4(n69), .Q(n789)
         );
  AO22X1 U813 ( .IN1(n2114), .IN2(n2226), .IN3(reg24[7]), .IN4(n69), .Q(n790)
         );
  AO22X1 U814 ( .IN1(n2115), .IN2(n2229), .IN3(reg24[8]), .IN4(n2113), .Q(n791) );
  AO22X1 U815 ( .IN1(n2115), .IN2(n2232), .IN3(reg24[9]), .IN4(n2113), .Q(n792) );
  AO22X1 U816 ( .IN1(n2114), .IN2(n2235), .IN3(reg24[10]), .IN4(n2113), .Q(
        n793) );
  AO22X1 U817 ( .IN1(n2114), .IN2(n2238), .IN3(reg24[11]), .IN4(n2113), .Q(
        n794) );
  AO22X1 U818 ( .IN1(n2114), .IN2(n2241), .IN3(reg24[12]), .IN4(n2113), .Q(
        n795) );
  AO22X1 U819 ( .IN1(n2114), .IN2(n2244), .IN3(reg24[13]), .IN4(n2113), .Q(
        n796) );
  AO22X1 U820 ( .IN1(n2114), .IN2(n2247), .IN3(reg24[14]), .IN4(n2113), .Q(
        n797) );
  AO22X1 U821 ( .IN1(n2114), .IN2(n2250), .IN3(reg24[15]), .IN4(n2113), .Q(
        n798) );
  AO22X1 U822 ( .IN1(n2114), .IN2(n2253), .IN3(reg24[16]), .IN4(n2113), .Q(
        n799) );
  AO22X1 U823 ( .IN1(n2114), .IN2(n2256), .IN3(reg24[17]), .IN4(n2113), .Q(
        n800) );
  AO22X1 U824 ( .IN1(n2114), .IN2(n2259), .IN3(reg24[18]), .IN4(n2113), .Q(
        n801) );
  AO22X1 U825 ( .IN1(n2115), .IN2(n2262), .IN3(reg24[19]), .IN4(n2113), .Q(
        n802) );
  AO22X1 U826 ( .IN1(n2114), .IN2(n2265), .IN3(reg24[20]), .IN4(n2112), .Q(
        n803) );
  AO22X1 U827 ( .IN1(n2115), .IN2(n2268), .IN3(reg24[21]), .IN4(n2112), .Q(
        n804) );
  AO22X1 U828 ( .IN1(n2114), .IN2(n2271), .IN3(reg24[22]), .IN4(n2112), .Q(
        n805) );
  AO22X1 U829 ( .IN1(n2115), .IN2(n2274), .IN3(reg24[23]), .IN4(n2112), .Q(
        n806) );
  AO22X1 U830 ( .IN1(n2114), .IN2(n2277), .IN3(reg24[24]), .IN4(n2112), .Q(
        n807) );
  AO22X1 U831 ( .IN1(n2115), .IN2(n2280), .IN3(reg24[25]), .IN4(n2112), .Q(
        n808) );
  AO22X1 U832 ( .IN1(n2115), .IN2(n2283), .IN3(reg24[26]), .IN4(n2112), .Q(
        n809) );
  AO22X1 U833 ( .IN1(n2115), .IN2(n2286), .IN3(reg24[27]), .IN4(n2112), .Q(
        n810) );
  AO22X1 U834 ( .IN1(n2115), .IN2(n2289), .IN3(reg24[28]), .IN4(n2112), .Q(
        n811) );
  AO22X1 U835 ( .IN1(n2115), .IN2(n2292), .IN3(reg24[29]), .IN4(n2112), .Q(
        n812) );
  AO22X1 U836 ( .IN1(n2115), .IN2(n2295), .IN3(reg24[30]), .IN4(n2112), .Q(
        n813) );
  AO22X1 U837 ( .IN1(n2115), .IN2(n2298), .IN3(reg24[31]), .IN4(n2112), .Q(
        n814) );
  AND3X1 U838 ( .IN1(wr_en), .IN2(n2392), .IN3(wr_addr[4]), .Q(n62) );
  AO22X1 U839 ( .IN1(n2111), .IN2(n2205), .IN3(reg25[0]), .IN4(n70), .Q(n815)
         );
  AO22X1 U840 ( .IN1(n2110), .IN2(n2208), .IN3(reg25[1]), .IN4(n70), .Q(n816)
         );
  AO22X1 U841 ( .IN1(n2111), .IN2(n2211), .IN3(reg25[2]), .IN4(n70), .Q(n817)
         );
  AO22X1 U842 ( .IN1(n2110), .IN2(n2214), .IN3(reg25[3]), .IN4(n70), .Q(n818)
         );
  AO22X1 U843 ( .IN1(n2110), .IN2(n2217), .IN3(reg25[4]), .IN4(n70), .Q(n819)
         );
  AO22X1 U844 ( .IN1(n2111), .IN2(n2220), .IN3(reg25[5]), .IN4(n70), .Q(n820)
         );
  AO22X1 U845 ( .IN1(n2111), .IN2(n2223), .IN3(reg25[6]), .IN4(n70), .Q(n821)
         );
  AO22X1 U846 ( .IN1(n2110), .IN2(n2226), .IN3(reg25[7]), .IN4(n70), .Q(n822)
         );
  AO22X1 U847 ( .IN1(n2111), .IN2(n2229), .IN3(reg25[8]), .IN4(n2109), .Q(n823) );
  AO22X1 U848 ( .IN1(n2111), .IN2(n2232), .IN3(reg25[9]), .IN4(n2109), .Q(n824) );
  AO22X1 U849 ( .IN1(n2110), .IN2(n2235), .IN3(reg25[10]), .IN4(n2109), .Q(
        n825) );
  AO22X1 U850 ( .IN1(n2110), .IN2(n2238), .IN3(reg25[11]), .IN4(n2109), .Q(
        n826) );
  AO22X1 U851 ( .IN1(n2110), .IN2(n2241), .IN3(reg25[12]), .IN4(n2109), .Q(
        n827) );
  AO22X1 U852 ( .IN1(n2110), .IN2(n2244), .IN3(reg25[13]), .IN4(n2109), .Q(
        n828) );
  AO22X1 U853 ( .IN1(n2110), .IN2(n2247), .IN3(reg25[14]), .IN4(n2109), .Q(
        n829) );
  AO22X1 U854 ( .IN1(n2110), .IN2(n2250), .IN3(reg25[15]), .IN4(n2109), .Q(
        n830) );
  AO22X1 U855 ( .IN1(n2110), .IN2(n2253), .IN3(reg25[16]), .IN4(n2109), .Q(
        n831) );
  AO22X1 U856 ( .IN1(n2110), .IN2(n2256), .IN3(reg25[17]), .IN4(n2109), .Q(
        n832) );
  AO22X1 U857 ( .IN1(n2110), .IN2(n2259), .IN3(reg25[18]), .IN4(n2109), .Q(
        n833) );
  AO22X1 U858 ( .IN1(n2111), .IN2(n2262), .IN3(reg25[19]), .IN4(n2109), .Q(
        n834) );
  AO22X1 U859 ( .IN1(n2110), .IN2(n2265), .IN3(reg25[20]), .IN4(n2108), .Q(
        n835) );
  AO22X1 U860 ( .IN1(n2111), .IN2(n2268), .IN3(reg25[21]), .IN4(n2108), .Q(
        n836) );
  AO22X1 U861 ( .IN1(n2110), .IN2(n2271), .IN3(reg25[22]), .IN4(n2108), .Q(
        n837) );
  AO22X1 U862 ( .IN1(n2111), .IN2(n2274), .IN3(reg25[23]), .IN4(n2108), .Q(
        n838) );
  AO22X1 U863 ( .IN1(n2110), .IN2(n2277), .IN3(reg25[24]), .IN4(n2108), .Q(
        n839) );
  AO22X1 U864 ( .IN1(n2111), .IN2(n2280), .IN3(reg25[25]), .IN4(n2108), .Q(
        n840) );
  AO22X1 U865 ( .IN1(n2111), .IN2(n2283), .IN3(reg25[26]), .IN4(n2108), .Q(
        n841) );
  AO22X1 U866 ( .IN1(n2111), .IN2(n2286), .IN3(reg25[27]), .IN4(n2108), .Q(
        n842) );
  AO22X1 U867 ( .IN1(n2111), .IN2(n2289), .IN3(reg25[28]), .IN4(n2108), .Q(
        n843) );
  AO22X1 U868 ( .IN1(n2111), .IN2(n2292), .IN3(reg25[29]), .IN4(n2108), .Q(
        n844) );
  AO22X1 U869 ( .IN1(n2111), .IN2(n2295), .IN3(reg25[30]), .IN4(n2108), .Q(
        n845) );
  AO22X1 U870 ( .IN1(n2111), .IN2(n2298), .IN3(reg25[31]), .IN4(n2108), .Q(
        n846) );
  NOR3X0 U871 ( .IN1(wr_addr[1]), .IN2(wr_addr[2]), .IN3(wr_addr[0]), .QN(n36)
         );
  AO22X1 U872 ( .IN1(n2107), .IN2(n2206), .IN3(reg26[0]), .IN4(n72), .Q(n847)
         );
  AO22X1 U873 ( .IN1(n2106), .IN2(n2209), .IN3(reg26[1]), .IN4(n72), .Q(n848)
         );
  AO22X1 U874 ( .IN1(n2107), .IN2(n2212), .IN3(reg26[2]), .IN4(n72), .Q(n849)
         );
  AO22X1 U875 ( .IN1(n2106), .IN2(n2215), .IN3(reg26[3]), .IN4(n72), .Q(n850)
         );
  AO22X1 U876 ( .IN1(n2106), .IN2(n2218), .IN3(reg26[4]), .IN4(n72), .Q(n851)
         );
  AO22X1 U877 ( .IN1(n2107), .IN2(n2221), .IN3(reg26[5]), .IN4(n72), .Q(n852)
         );
  AO22X1 U878 ( .IN1(n2107), .IN2(n2224), .IN3(reg26[6]), .IN4(n72), .Q(n853)
         );
  AO22X1 U879 ( .IN1(n2106), .IN2(n2227), .IN3(reg26[7]), .IN4(n72), .Q(n854)
         );
  AO22X1 U880 ( .IN1(n2107), .IN2(n2230), .IN3(reg26[8]), .IN4(n2105), .Q(n855) );
  AO22X1 U881 ( .IN1(n2107), .IN2(n2233), .IN3(reg26[9]), .IN4(n2105), .Q(n856) );
  AO22X1 U882 ( .IN1(n2106), .IN2(n2236), .IN3(reg26[10]), .IN4(n2105), .Q(
        n857) );
  AO22X1 U883 ( .IN1(n2106), .IN2(n2239), .IN3(reg26[11]), .IN4(n2105), .Q(
        n858) );
  AO22X1 U884 ( .IN1(n2106), .IN2(n2242), .IN3(reg26[12]), .IN4(n2105), .Q(
        n859) );
  AO22X1 U885 ( .IN1(n2106), .IN2(n2245), .IN3(reg26[13]), .IN4(n2105), .Q(
        n860) );
  AO22X1 U886 ( .IN1(n2106), .IN2(n2248), .IN3(reg26[14]), .IN4(n2105), .Q(
        n861) );
  AO22X1 U887 ( .IN1(n2106), .IN2(n2251), .IN3(reg26[15]), .IN4(n2105), .Q(
        n862) );
  AO22X1 U888 ( .IN1(n2106), .IN2(n2254), .IN3(reg26[16]), .IN4(n2105), .Q(
        n863) );
  AO22X1 U889 ( .IN1(n2106), .IN2(n2257), .IN3(reg26[17]), .IN4(n2105), .Q(
        n864) );
  AO22X1 U890 ( .IN1(n2106), .IN2(n2260), .IN3(reg26[18]), .IN4(n2105), .Q(
        n865) );
  AO22X1 U891 ( .IN1(n2107), .IN2(n2263), .IN3(reg26[19]), .IN4(n2105), .Q(
        n866) );
  AO22X1 U892 ( .IN1(n2106), .IN2(n2266), .IN3(reg26[20]), .IN4(n2104), .Q(
        n867) );
  AO22X1 U893 ( .IN1(n2107), .IN2(n2269), .IN3(reg26[21]), .IN4(n2104), .Q(
        n868) );
  AO22X1 U894 ( .IN1(n2106), .IN2(n2272), .IN3(reg26[22]), .IN4(n2104), .Q(
        n869) );
  AO22X1 U895 ( .IN1(n2107), .IN2(n2275), .IN3(reg26[23]), .IN4(n2104), .Q(
        n870) );
  AO22X1 U896 ( .IN1(n2106), .IN2(n2278), .IN3(reg26[24]), .IN4(n2104), .Q(
        n871) );
  AO22X1 U897 ( .IN1(n2107), .IN2(n2281), .IN3(reg26[25]), .IN4(n2104), .Q(
        n872) );
  AO22X1 U898 ( .IN1(n2107), .IN2(n2284), .IN3(reg26[26]), .IN4(n2104), .Q(
        n873) );
  AO22X1 U899 ( .IN1(n2107), .IN2(n2287), .IN3(reg26[27]), .IN4(n2104), .Q(
        n874) );
  AO22X1 U900 ( .IN1(n2107), .IN2(n2290), .IN3(reg26[28]), .IN4(n2104), .Q(
        n875) );
  AO22X1 U901 ( .IN1(n2107), .IN2(n2293), .IN3(reg26[29]), .IN4(n2104), .Q(
        n876) );
  AO22X1 U902 ( .IN1(n2107), .IN2(n2296), .IN3(reg26[30]), .IN4(n2104), .Q(
        n877) );
  AO22X1 U903 ( .IN1(n2107), .IN2(n2299), .IN3(reg26[31]), .IN4(n2104), .Q(
        n878) );
  NOR3X0 U904 ( .IN1(wr_addr[1]), .IN2(wr_addr[2]), .IN3(n2390), .QN(n38) );
  AO22X1 U905 ( .IN1(n2103), .IN2(n2206), .IN3(reg27[0]), .IN4(n73), .Q(n879)
         );
  AO22X1 U906 ( .IN1(n2102), .IN2(n2209), .IN3(reg27[1]), .IN4(n73), .Q(n880)
         );
  AO22X1 U907 ( .IN1(n2103), .IN2(n2212), .IN3(reg27[2]), .IN4(n73), .Q(n881)
         );
  AO22X1 U908 ( .IN1(n2102), .IN2(n2215), .IN3(reg27[3]), .IN4(n73), .Q(n882)
         );
  AO22X1 U909 ( .IN1(n2102), .IN2(n2218), .IN3(reg27[4]), .IN4(n73), .Q(n883)
         );
  AO22X1 U910 ( .IN1(n2103), .IN2(n2221), .IN3(reg27[5]), .IN4(n73), .Q(n884)
         );
  AO22X1 U911 ( .IN1(n2103), .IN2(n2224), .IN3(reg27[6]), .IN4(n73), .Q(n885)
         );
  AO22X1 U912 ( .IN1(n2102), .IN2(n2227), .IN3(reg27[7]), .IN4(n73), .Q(n886)
         );
  AO22X1 U913 ( .IN1(n2103), .IN2(n2230), .IN3(reg27[8]), .IN4(n2101), .Q(n887) );
  AO22X1 U914 ( .IN1(n2103), .IN2(n2233), .IN3(reg27[9]), .IN4(n2101), .Q(n888) );
  AO22X1 U915 ( .IN1(n2102), .IN2(n2236), .IN3(reg27[10]), .IN4(n2101), .Q(
        n889) );
  AO22X1 U916 ( .IN1(n2102), .IN2(n2239), .IN3(reg27[11]), .IN4(n2101), .Q(
        n890) );
  AO22X1 U917 ( .IN1(n2102), .IN2(n2242), .IN3(reg27[12]), .IN4(n2101), .Q(
        n891) );
  AO22X1 U918 ( .IN1(n2102), .IN2(n2245), .IN3(reg27[13]), .IN4(n2101), .Q(
        n892) );
  AO22X1 U919 ( .IN1(n2102), .IN2(n2248), .IN3(reg27[14]), .IN4(n2101), .Q(
        n893) );
  AO22X1 U920 ( .IN1(n2102), .IN2(n2251), .IN3(reg27[15]), .IN4(n2101), .Q(
        n894) );
  AO22X1 U921 ( .IN1(n2102), .IN2(n2254), .IN3(reg27[16]), .IN4(n2101), .Q(
        n895) );
  AO22X1 U922 ( .IN1(n2102), .IN2(n2257), .IN3(reg27[17]), .IN4(n2101), .Q(
        n896) );
  AO22X1 U923 ( .IN1(n2102), .IN2(n2260), .IN3(reg27[18]), .IN4(n2101), .Q(
        n897) );
  AO22X1 U924 ( .IN1(n2103), .IN2(n2263), .IN3(reg27[19]), .IN4(n2101), .Q(
        n898) );
  AO22X1 U925 ( .IN1(n2102), .IN2(n2266), .IN3(reg27[20]), .IN4(n2100), .Q(
        n899) );
  AO22X1 U926 ( .IN1(n2103), .IN2(n2269), .IN3(reg27[21]), .IN4(n2100), .Q(
        n900) );
  AO22X1 U927 ( .IN1(n2102), .IN2(n2272), .IN3(reg27[22]), .IN4(n2100), .Q(
        n901) );
  AO22X1 U928 ( .IN1(n2103), .IN2(n2275), .IN3(reg27[23]), .IN4(n2100), .Q(
        n902) );
  AO22X1 U929 ( .IN1(n2102), .IN2(n2278), .IN3(reg27[24]), .IN4(n2100), .Q(
        n903) );
  AO22X1 U930 ( .IN1(n2103), .IN2(n2281), .IN3(reg27[25]), .IN4(n2100), .Q(
        n904) );
  AO22X1 U931 ( .IN1(n2103), .IN2(n2284), .IN3(reg27[26]), .IN4(n2100), .Q(
        n905) );
  AO22X1 U932 ( .IN1(n2103), .IN2(n2287), .IN3(reg27[27]), .IN4(n2100), .Q(
        n906) );
  AO22X1 U933 ( .IN1(n2103), .IN2(n2290), .IN3(reg27[28]), .IN4(n2100), .Q(
        n907) );
  AO22X1 U934 ( .IN1(n2103), .IN2(n2293), .IN3(reg27[29]), .IN4(n2100), .Q(
        n908) );
  AO22X1 U935 ( .IN1(n2103), .IN2(n2296), .IN3(reg27[30]), .IN4(n2100), .Q(
        n909) );
  AO22X1 U936 ( .IN1(n2103), .IN2(n2299), .IN3(reg27[31]), .IN4(n2100), .Q(
        n910) );
  NOR3X0 U937 ( .IN1(wr_addr[0]), .IN2(wr_addr[2]), .IN3(n2391), .QN(n41) );
  AO22X1 U938 ( .IN1(n2099), .IN2(n2206), .IN3(reg28[0]), .IN4(n74), .Q(n911)
         );
  AO22X1 U939 ( .IN1(n2098), .IN2(n2209), .IN3(reg28[1]), .IN4(n74), .Q(n912)
         );
  AO22X1 U940 ( .IN1(n2099), .IN2(n2212), .IN3(reg28[2]), .IN4(n74), .Q(n913)
         );
  AO22X1 U941 ( .IN1(n2098), .IN2(n2215), .IN3(reg28[3]), .IN4(n74), .Q(n914)
         );
  AO22X1 U942 ( .IN1(n2098), .IN2(n2218), .IN3(reg28[4]), .IN4(n74), .Q(n915)
         );
  AO22X1 U943 ( .IN1(n2099), .IN2(n2221), .IN3(reg28[5]), .IN4(n74), .Q(n916)
         );
  AO22X1 U944 ( .IN1(n2099), .IN2(n2224), .IN3(reg28[6]), .IN4(n74), .Q(n917)
         );
  AO22X1 U945 ( .IN1(n2098), .IN2(n2227), .IN3(reg28[7]), .IN4(n74), .Q(n918)
         );
  AO22X1 U946 ( .IN1(n2099), .IN2(n2230), .IN3(reg28[8]), .IN4(n2097), .Q(n919) );
  AO22X1 U947 ( .IN1(n2099), .IN2(n2233), .IN3(reg28[9]), .IN4(n2097), .Q(n920) );
  AO22X1 U948 ( .IN1(n2098), .IN2(n2236), .IN3(reg28[10]), .IN4(n2097), .Q(
        n921) );
  AO22X1 U949 ( .IN1(n2098), .IN2(n2239), .IN3(reg28[11]), .IN4(n2097), .Q(
        n922) );
  AO22X1 U950 ( .IN1(n2098), .IN2(n2242), .IN3(reg28[12]), .IN4(n2097), .Q(
        n923) );
  AO22X1 U951 ( .IN1(n2098), .IN2(n2245), .IN3(reg28[13]), .IN4(n2097), .Q(
        n924) );
  AO22X1 U952 ( .IN1(n2098), .IN2(n2248), .IN3(reg28[14]), .IN4(n2097), .Q(
        n925) );
  AO22X1 U953 ( .IN1(n2098), .IN2(n2251), .IN3(reg28[15]), .IN4(n2097), .Q(
        n926) );
  AO22X1 U954 ( .IN1(n2098), .IN2(n2254), .IN3(reg28[16]), .IN4(n2097), .Q(
        n927) );
  AO22X1 U955 ( .IN1(n2098), .IN2(n2257), .IN3(reg28[17]), .IN4(n2097), .Q(
        n928) );
  AO22X1 U956 ( .IN1(n2098), .IN2(n2260), .IN3(reg28[18]), .IN4(n2097), .Q(
        n929) );
  AO22X1 U957 ( .IN1(n2099), .IN2(n2263), .IN3(reg28[19]), .IN4(n2097), .Q(
        n930) );
  AO22X1 U958 ( .IN1(n2098), .IN2(n2266), .IN3(reg28[20]), .IN4(n2096), .Q(
        n931) );
  AO22X1 U959 ( .IN1(n2099), .IN2(n2269), .IN3(reg28[21]), .IN4(n2096), .Q(
        n932) );
  AO22X1 U960 ( .IN1(n2098), .IN2(n2272), .IN3(reg28[22]), .IN4(n2096), .Q(
        n933) );
  AO22X1 U961 ( .IN1(n2099), .IN2(n2275), .IN3(reg28[23]), .IN4(n2096), .Q(
        n934) );
  AO22X1 U962 ( .IN1(n2098), .IN2(n2278), .IN3(reg28[24]), .IN4(n2096), .Q(
        n935) );
  AO22X1 U963 ( .IN1(n2099), .IN2(n2281), .IN3(reg28[25]), .IN4(n2096), .Q(
        n936) );
  AO22X1 U964 ( .IN1(n2099), .IN2(n2284), .IN3(reg28[26]), .IN4(n2096), .Q(
        n937) );
  AO22X1 U965 ( .IN1(n2099), .IN2(n2287), .IN3(reg28[27]), .IN4(n2096), .Q(
        n938) );
  AO22X1 U966 ( .IN1(n2099), .IN2(n2290), .IN3(reg28[28]), .IN4(n2096), .Q(
        n939) );
  AO22X1 U967 ( .IN1(n2099), .IN2(n2293), .IN3(reg28[29]), .IN4(n2096), .Q(
        n940) );
  AO22X1 U968 ( .IN1(n2099), .IN2(n2296), .IN3(reg28[30]), .IN4(n2096), .Q(
        n941) );
  AO22X1 U969 ( .IN1(n2099), .IN2(n2299), .IN3(reg28[31]), .IN4(n2096), .Q(
        n942) );
  NOR3X0 U970 ( .IN1(n2390), .IN2(wr_addr[2]), .IN3(n2391), .QN(n43) );
  AO22X1 U971 ( .IN1(n2095), .IN2(n2206), .IN3(reg29[0]), .IN4(n75), .Q(n943)
         );
  AO22X1 U972 ( .IN1(n2094), .IN2(n2209), .IN3(reg29[1]), .IN4(n75), .Q(n944)
         );
  AO22X1 U973 ( .IN1(n2095), .IN2(n2212), .IN3(reg29[2]), .IN4(n75), .Q(n945)
         );
  AO22X1 U974 ( .IN1(n2094), .IN2(n2215), .IN3(reg29[3]), .IN4(n75), .Q(n946)
         );
  AO22X1 U975 ( .IN1(n2094), .IN2(n2218), .IN3(reg29[4]), .IN4(n75), .Q(n947)
         );
  AO22X1 U976 ( .IN1(n2095), .IN2(n2221), .IN3(reg29[5]), .IN4(n75), .Q(n948)
         );
  AO22X1 U977 ( .IN1(n2095), .IN2(n2224), .IN3(reg29[6]), .IN4(n75), .Q(n949)
         );
  AO22X1 U978 ( .IN1(n2094), .IN2(n2227), .IN3(reg29[7]), .IN4(n75), .Q(n950)
         );
  AO22X1 U979 ( .IN1(n2095), .IN2(n2230), .IN3(reg29[8]), .IN4(n2093), .Q(n951) );
  AO22X1 U980 ( .IN1(n2095), .IN2(n2233), .IN3(reg29[9]), .IN4(n2093), .Q(n952) );
  AO22X1 U981 ( .IN1(n2094), .IN2(n2236), .IN3(reg29[10]), .IN4(n2093), .Q(
        n953) );
  AO22X1 U982 ( .IN1(n2094), .IN2(n2239), .IN3(reg29[11]), .IN4(n2093), .Q(
        n954) );
  AO22X1 U983 ( .IN1(n2094), .IN2(n2242), .IN3(reg29[12]), .IN4(n2093), .Q(
        n955) );
  AO22X1 U984 ( .IN1(n2094), .IN2(n2245), .IN3(reg29[13]), .IN4(n2093), .Q(
        n956) );
  AO22X1 U985 ( .IN1(n2094), .IN2(n2248), .IN3(reg29[14]), .IN4(n2093), .Q(
        n957) );
  AO22X1 U986 ( .IN1(n2094), .IN2(n2251), .IN3(reg29[15]), .IN4(n2093), .Q(
        n958) );
  AO22X1 U987 ( .IN1(n2094), .IN2(n2254), .IN3(reg29[16]), .IN4(n2093), .Q(
        n959) );
  AO22X1 U988 ( .IN1(n2094), .IN2(n2257), .IN3(reg29[17]), .IN4(n2093), .Q(
        n960) );
  AO22X1 U989 ( .IN1(n2094), .IN2(n2260), .IN3(reg29[18]), .IN4(n2093), .Q(
        n961) );
  AO22X1 U990 ( .IN1(n2095), .IN2(n2263), .IN3(reg29[19]), .IN4(n2093), .Q(
        n962) );
  AO22X1 U991 ( .IN1(n2094), .IN2(n2266), .IN3(reg29[20]), .IN4(n2092), .Q(
        n963) );
  AO22X1 U992 ( .IN1(n2095), .IN2(n2269), .IN3(reg29[21]), .IN4(n2092), .Q(
        n964) );
  AO22X1 U993 ( .IN1(n2094), .IN2(n2272), .IN3(reg29[22]), .IN4(n2092), .Q(
        n965) );
  AO22X1 U994 ( .IN1(n2095), .IN2(n2275), .IN3(reg29[23]), .IN4(n2092), .Q(
        n966) );
  AO22X1 U995 ( .IN1(n2094), .IN2(n2278), .IN3(reg29[24]), .IN4(n2092), .Q(
        n967) );
  AO22X1 U996 ( .IN1(n2095), .IN2(n2281), .IN3(reg29[25]), .IN4(n2092), .Q(
        n968) );
  AO22X1 U997 ( .IN1(n2095), .IN2(n2284), .IN3(reg29[26]), .IN4(n2092), .Q(
        n969) );
  AO22X1 U998 ( .IN1(n2095), .IN2(n2287), .IN3(reg29[27]), .IN4(n2092), .Q(
        n970) );
  AO22X1 U999 ( .IN1(n2095), .IN2(n2290), .IN3(reg29[28]), .IN4(n2092), .Q(
        n971) );
  AO22X1 U1000 ( .IN1(n2095), .IN2(n2293), .IN3(reg29[29]), .IN4(n2092), .Q(
        n972) );
  AO22X1 U1001 ( .IN1(n2095), .IN2(n2296), .IN3(reg29[30]), .IN4(n2092), .Q(
        n973) );
  AO22X1 U1002 ( .IN1(n2095), .IN2(n2299), .IN3(reg29[31]), .IN4(n2092), .Q(
        n974) );
  AND3X1 U1003 ( .IN1(n2390), .IN2(n2391), .IN3(wr_addr[2]), .Q(n45) );
  AO22X1 U1004 ( .IN1(n2091), .IN2(n2206), .IN3(reg30[0]), .IN4(n76), .Q(n975)
         );
  AO22X1 U1005 ( .IN1(n2090), .IN2(n2209), .IN3(reg30[1]), .IN4(n76), .Q(n976)
         );
  AO22X1 U1006 ( .IN1(n2091), .IN2(n2212), .IN3(reg30[2]), .IN4(n76), .Q(n977)
         );
  AO22X1 U1007 ( .IN1(n2090), .IN2(n2215), .IN3(reg30[3]), .IN4(n76), .Q(n978)
         );
  AO22X1 U1008 ( .IN1(n2090), .IN2(n2218), .IN3(reg30[4]), .IN4(n76), .Q(n979)
         );
  AO22X1 U1009 ( .IN1(n2091), .IN2(n2221), .IN3(reg30[5]), .IN4(n76), .Q(n980)
         );
  AO22X1 U1010 ( .IN1(n2091), .IN2(n2224), .IN3(reg30[6]), .IN4(n76), .Q(n981)
         );
  AO22X1 U1011 ( .IN1(n2090), .IN2(n2227), .IN3(reg30[7]), .IN4(n76), .Q(n982)
         );
  AO22X1 U1012 ( .IN1(n2091), .IN2(n2230), .IN3(reg30[8]), .IN4(n2089), .Q(
        n983) );
  AO22X1 U1013 ( .IN1(n2091), .IN2(n2233), .IN3(reg30[9]), .IN4(n2089), .Q(
        n984) );
  AO22X1 U1014 ( .IN1(n2090), .IN2(n2236), .IN3(reg30[10]), .IN4(n2089), .Q(
        n985) );
  AO22X1 U1015 ( .IN1(n2090), .IN2(n2239), .IN3(reg30[11]), .IN4(n2089), .Q(
        n986) );
  AO22X1 U1016 ( .IN1(n2090), .IN2(n2242), .IN3(reg30[12]), .IN4(n2089), .Q(
        n987) );
  AO22X1 U1017 ( .IN1(n2090), .IN2(n2245), .IN3(reg30[13]), .IN4(n2089), .Q(
        n988) );
  AO22X1 U1018 ( .IN1(n2090), .IN2(n2248), .IN3(reg30[14]), .IN4(n2089), .Q(
        n989) );
  AO22X1 U1019 ( .IN1(n2090), .IN2(n2251), .IN3(reg30[15]), .IN4(n2089), .Q(
        n990) );
  AO22X1 U1020 ( .IN1(n2090), .IN2(n2254), .IN3(reg30[16]), .IN4(n2089), .Q(
        n991) );
  AO22X1 U1021 ( .IN1(n2090), .IN2(n2257), .IN3(reg30[17]), .IN4(n2089), .Q(
        n992) );
  AO22X1 U1022 ( .IN1(n2090), .IN2(n2260), .IN3(reg30[18]), .IN4(n2089), .Q(
        n993) );
  AO22X1 U1023 ( .IN1(n2091), .IN2(n2263), .IN3(reg30[19]), .IN4(n2089), .Q(
        n994) );
  AO22X1 U1024 ( .IN1(n2090), .IN2(n2266), .IN3(reg30[20]), .IN4(n2088), .Q(
        n995) );
  AO22X1 U1025 ( .IN1(n2091), .IN2(n2269), .IN3(reg30[21]), .IN4(n2088), .Q(
        n996) );
  AO22X1 U1026 ( .IN1(n2090), .IN2(n2272), .IN3(reg30[22]), .IN4(n2088), .Q(
        n997) );
  AO22X1 U1027 ( .IN1(n2091), .IN2(n2275), .IN3(reg30[23]), .IN4(n2088), .Q(
        n998) );
  AO22X1 U1028 ( .IN1(n2090), .IN2(n2278), .IN3(reg30[24]), .IN4(n2088), .Q(
        n999) );
  AO22X1 U1029 ( .IN1(n2091), .IN2(n2281), .IN3(reg30[25]), .IN4(n2088), .Q(
        n1000) );
  AO22X1 U1030 ( .IN1(n2091), .IN2(n2284), .IN3(reg30[26]), .IN4(n2088), .Q(
        n1001) );
  AO22X1 U1031 ( .IN1(n2091), .IN2(n2287), .IN3(reg30[27]), .IN4(n2088), .Q(
        n1002) );
  AO22X1 U1032 ( .IN1(n2091), .IN2(n2290), .IN3(reg30[28]), .IN4(n2088), .Q(
        n1003) );
  AO22X1 U1033 ( .IN1(n2091), .IN2(n2293), .IN3(reg30[29]), .IN4(n2088), .Q(
        n1004) );
  AO22X1 U1034 ( .IN1(n2091), .IN2(n2296), .IN3(reg30[30]), .IN4(n2088), .Q(
        n1005) );
  AO22X1 U1035 ( .IN1(n2091), .IN2(n2299), .IN3(reg30[31]), .IN4(n2088), .Q(
        n1006) );
  AND3X1 U1036 ( .IN1(wr_addr[0]), .IN2(n2391), .IN3(wr_addr[2]), .Q(n47) );
  AO22X1 U1037 ( .IN1(n2087), .IN2(n2206), .IN3(reg31[0]), .IN4(n77), .Q(n1007) );
  AO22X1 U1038 ( .IN1(n2086), .IN2(n2209), .IN3(reg31[1]), .IN4(n77), .Q(n1008) );
  AO22X1 U1039 ( .IN1(n2087), .IN2(n2212), .IN3(reg31[2]), .IN4(n77), .Q(n1009) );
  AO22X1 U1040 ( .IN1(n2086), .IN2(n2215), .IN3(reg31[3]), .IN4(n77), .Q(n1010) );
  AO22X1 U1041 ( .IN1(n2086), .IN2(n2218), .IN3(reg31[4]), .IN4(n77), .Q(n1011) );
  AO22X1 U1042 ( .IN1(n2087), .IN2(n2221), .IN3(reg31[5]), .IN4(n77), .Q(n1012) );
  AO22X1 U1043 ( .IN1(n2087), .IN2(n2224), .IN3(reg31[6]), .IN4(n77), .Q(n1013) );
  AO22X1 U1044 ( .IN1(n2086), .IN2(n2227), .IN3(reg31[7]), .IN4(n77), .Q(n1014) );
  AO22X1 U1045 ( .IN1(n2087), .IN2(n2230), .IN3(reg31[8]), .IN4(n2085), .Q(
        n1015) );
  AO22X1 U1046 ( .IN1(n2087), .IN2(n2233), .IN3(reg31[9]), .IN4(n2085), .Q(
        n1016) );
  AO22X1 U1047 ( .IN1(n2086), .IN2(n2236), .IN3(reg31[10]), .IN4(n2085), .Q(
        n1017) );
  AO22X1 U1048 ( .IN1(n2086), .IN2(n2239), .IN3(reg31[11]), .IN4(n2085), .Q(
        n1018) );
  AO22X1 U1049 ( .IN1(n2086), .IN2(n2242), .IN3(reg31[12]), .IN4(n2085), .Q(
        n1019) );
  AO22X1 U1050 ( .IN1(n2086), .IN2(n2245), .IN3(reg31[13]), .IN4(n2085), .Q(
        n1020) );
  AO22X1 U1051 ( .IN1(n2086), .IN2(n2248), .IN3(reg31[14]), .IN4(n2085), .Q(
        n1021) );
  AO22X1 U1052 ( .IN1(n2086), .IN2(n2251), .IN3(reg31[15]), .IN4(n2085), .Q(
        n1022) );
  AO22X1 U1053 ( .IN1(n2086), .IN2(n2254), .IN3(reg31[16]), .IN4(n2085), .Q(
        n1023) );
  AO22X1 U1054 ( .IN1(n2086), .IN2(n2257), .IN3(reg31[17]), .IN4(n2085), .Q(
        n1024) );
  AO22X1 U1055 ( .IN1(n2086), .IN2(n2260), .IN3(reg31[18]), .IN4(n2085), .Q(
        n1025) );
  AO22X1 U1056 ( .IN1(n2087), .IN2(n2263), .IN3(reg31[19]), .IN4(n2085), .Q(
        n1026) );
  AO22X1 U1057 ( .IN1(n2086), .IN2(n2266), .IN3(reg31[20]), .IN4(n2084), .Q(
        n1027) );
  AO22X1 U1058 ( .IN1(n2087), .IN2(n2269), .IN3(reg31[21]), .IN4(n2084), .Q(
        n1028) );
  AO22X1 U1059 ( .IN1(n2086), .IN2(n2272), .IN3(reg31[22]), .IN4(n2084), .Q(
        n1029) );
  AO22X1 U1060 ( .IN1(n2087), .IN2(n2275), .IN3(reg31[23]), .IN4(n2084), .Q(
        n1030) );
  AO22X1 U1061 ( .IN1(n2086), .IN2(n2278), .IN3(reg31[24]), .IN4(n2084), .Q(
        n1031) );
  AO22X1 U1062 ( .IN1(n2087), .IN2(n2281), .IN3(reg31[25]), .IN4(n2084), .Q(
        n1032) );
  AO22X1 U1063 ( .IN1(n2087), .IN2(n2284), .IN3(reg31[26]), .IN4(n2084), .Q(
        n1033) );
  AO22X1 U1064 ( .IN1(n2087), .IN2(n2287), .IN3(reg31[27]), .IN4(n2084), .Q(
        n1034) );
  AO22X1 U1065 ( .IN1(n2087), .IN2(n2290), .IN3(reg31[28]), .IN4(n2084), .Q(
        n1035) );
  AO22X1 U1066 ( .IN1(n2087), .IN2(n2293), .IN3(reg31[29]), .IN4(n2084), .Q(
        n1036) );
  AO22X1 U1067 ( .IN1(n2087), .IN2(n2296), .IN3(reg31[30]), .IN4(n2084), .Q(
        n1037) );
  AO22X1 U1068 ( .IN1(n2087), .IN2(n2299), .IN3(reg31[31]), .IN4(n2084), .Q(
        n1038) );
  AND3X1 U1069 ( .IN1(wr_addr[1]), .IN2(n2390), .IN3(wr_addr[2]), .Q(n49) );
  AO22X1 U1070 ( .IN1(n2083), .IN2(n2206), .IN3(reg32[0]), .IN4(n78), .Q(n1039) );
  AO22X1 U1071 ( .IN1(n2082), .IN2(n2209), .IN3(reg32[1]), .IN4(n78), .Q(n1040) );
  AO22X1 U1072 ( .IN1(n2083), .IN2(n2212), .IN3(reg32[2]), .IN4(n78), .Q(n1041) );
  AO22X1 U1073 ( .IN1(n2082), .IN2(n2215), .IN3(reg32[3]), .IN4(n78), .Q(n1042) );
  AO22X1 U1074 ( .IN1(n2082), .IN2(n2218), .IN3(reg32[4]), .IN4(n78), .Q(n1043) );
  AO22X1 U1075 ( .IN1(n2083), .IN2(n2221), .IN3(reg32[5]), .IN4(n78), .Q(n1044) );
  AO22X1 U1076 ( .IN1(n2083), .IN2(n2224), .IN3(reg32[6]), .IN4(n78), .Q(n1045) );
  AO22X1 U1077 ( .IN1(n2082), .IN2(n2227), .IN3(reg32[7]), .IN4(n78), .Q(n1046) );
  AO22X1 U1078 ( .IN1(n2083), .IN2(n2230), .IN3(reg32[8]), .IN4(n2081), .Q(
        n1047) );
  AO22X1 U1079 ( .IN1(n2083), .IN2(n2233), .IN3(reg32[9]), .IN4(n2081), .Q(
        n1048) );
  AO22X1 U1080 ( .IN1(n2082), .IN2(n2236), .IN3(reg32[10]), .IN4(n2081), .Q(
        n1049) );
  AO22X1 U1081 ( .IN1(n2082), .IN2(n2239), .IN3(reg32[11]), .IN4(n2081), .Q(
        n1050) );
  AO22X1 U1082 ( .IN1(n2082), .IN2(n2242), .IN3(reg32[12]), .IN4(n2081), .Q(
        n1051) );
  AO22X1 U1083 ( .IN1(n2082), .IN2(n2245), .IN3(reg32[13]), .IN4(n2081), .Q(
        n1052) );
  AO22X1 U1084 ( .IN1(n2082), .IN2(n2248), .IN3(reg32[14]), .IN4(n2081), .Q(
        n1053) );
  AO22X1 U1085 ( .IN1(n2082), .IN2(n2251), .IN3(reg32[15]), .IN4(n2081), .Q(
        n1054) );
  AO22X1 U1086 ( .IN1(n2082), .IN2(n2254), .IN3(reg32[16]), .IN4(n2081), .Q(
        n1055) );
  AO22X1 U1087 ( .IN1(n2082), .IN2(n2257), .IN3(reg32[17]), .IN4(n2081), .Q(
        n1056) );
  AO22X1 U1088 ( .IN1(n2082), .IN2(n2260), .IN3(reg32[18]), .IN4(n2081), .Q(
        n1057) );
  AO22X1 U1089 ( .IN1(n2083), .IN2(n2263), .IN3(reg32[19]), .IN4(n2081), .Q(
        n1058) );
  AO22X1 U1090 ( .IN1(n2082), .IN2(n2266), .IN3(reg32[20]), .IN4(n2080), .Q(
        n1059) );
  AO22X1 U1091 ( .IN1(n2083), .IN2(n2269), .IN3(reg32[21]), .IN4(n2080), .Q(
        n1060) );
  AO22X1 U1092 ( .IN1(n2082), .IN2(n2272), .IN3(reg32[22]), .IN4(n2080), .Q(
        n1061) );
  AO22X1 U1093 ( .IN1(n2083), .IN2(n2275), .IN3(reg32[23]), .IN4(n2080), .Q(
        n1062) );
  AO22X1 U1094 ( .IN1(n2082), .IN2(n2278), .IN3(reg32[24]), .IN4(n2080), .Q(
        n1063) );
  AO22X1 U1095 ( .IN1(n2083), .IN2(n2281), .IN3(reg32[25]), .IN4(n2080), .Q(
        n1064) );
  AO22X1 U1096 ( .IN1(n2083), .IN2(n2284), .IN3(reg32[26]), .IN4(n2080), .Q(
        n1065) );
  AO22X1 U1097 ( .IN1(n2083), .IN2(n2287), .IN3(reg32[27]), .IN4(n2080), .Q(
        n1066) );
  AO22X1 U1098 ( .IN1(n2083), .IN2(n2290), .IN3(reg32[28]), .IN4(n2080), .Q(
        n1067) );
  AO22X1 U1099 ( .IN1(n2083), .IN2(n2293), .IN3(reg32[29]), .IN4(n2080), .Q(
        n1068) );
  AO22X1 U1100 ( .IN1(n2083), .IN2(n2296), .IN3(reg32[30]), .IN4(n2080), .Q(
        n1069) );
  AO22X1 U1101 ( .IN1(n2083), .IN2(n2299), .IN3(reg32[31]), .IN4(n2080), .Q(
        n1070) );
  AND3X1 U1102 ( .IN1(wr_addr[1]), .IN2(wr_addr[0]), .IN3(wr_addr[2]), .Q(n51)
         );
  AND3X1 U1103 ( .IN1(wr_addr[3]), .IN2(wr_en), .IN3(wr_addr[4]), .Q(n71) );
  NAND2X0 U2 ( .IN1(n38), .IN2(n39), .QN(n37) );
  NAND2X0 U3 ( .IN1(n43), .IN2(n39), .QN(n42) );
  NAND2X0 U4 ( .IN1(n41), .IN2(n39), .QN(n40) );
  NAND2X0 U5 ( .IN1(n71), .IN2(n43), .QN(n74) );
  NAND2X0 U6 ( .IN1(n71), .IN2(n41), .QN(n73) );
  NAND2X0 U7 ( .IN1(n71), .IN2(n38), .QN(n72) );
  NAND2X0 U8 ( .IN1(n62), .IN2(n43), .QN(n65) );
  NAND2X0 U9 ( .IN1(n62), .IN2(n41), .QN(n64) );
  NAND2X0 U10 ( .IN1(n62), .IN2(n38), .QN(n63) );
  NAND2X0 U11 ( .IN1(n53), .IN2(n43), .QN(n56) );
  NAND2X0 U12 ( .IN1(n53), .IN2(n41), .QN(n55) );
  NAND2X0 U13 ( .IN1(n53), .IN2(n38), .QN(n54) );
  NAND2X0 U14 ( .IN1(n62), .IN2(n51), .QN(n69) );
  NAND2X0 U15 ( .IN1(n62), .IN2(n49), .QN(n68) );
  NAND2X0 U16 ( .IN1(n62), .IN2(n47), .QN(n67) );
  NAND2X0 U17 ( .IN1(n62), .IN2(n45), .QN(n66) );
  NAND2X0 U18 ( .IN1(n62), .IN2(n36), .QN(n61) );
  NAND2X0 U19 ( .IN1(n53), .IN2(n51), .QN(n60) );
  NAND2X0 U20 ( .IN1(n53), .IN2(n49), .QN(n59) );
  NAND2X0 U21 ( .IN1(n53), .IN2(n47), .QN(n58) );
  NAND2X0 U22 ( .IN1(n53), .IN2(n45), .QN(n57) );
  NAND2X0 U23 ( .IN1(n53), .IN2(n36), .QN(n52) );
  NAND2X0 U24 ( .IN1(n71), .IN2(n51), .QN(n78) );
  NAND2X0 U25 ( .IN1(n71), .IN2(n49), .QN(n77) );
  NAND2X0 U26 ( .IN1(n71), .IN2(n47), .QN(n76) );
  NAND2X0 U27 ( .IN1(n71), .IN2(n45), .QN(n75) );
  NAND2X0 U28 ( .IN1(n71), .IN2(n36), .QN(n70) );
  NAND2X0 U29 ( .IN1(n51), .IN2(n39), .QN(n50) );
  NAND2X0 U30 ( .IN1(n49), .IN2(n39), .QN(n48) );
  NAND2X0 U31 ( .IN1(n47), .IN2(n39), .QN(n46) );
  NAND2X0 U32 ( .IN1(n45), .IN2(n39), .QN(n44) );
  INVX0 U33 ( .INP(n37), .ZN(n2202) );
  INVX0 U34 ( .INP(n37), .ZN(n2203) );
  INVX0 U35 ( .INP(n40), .ZN(n2198) );
  INVX0 U36 ( .INP(n40), .ZN(n2199) );
  INVX0 U37 ( .INP(n42), .ZN(n2194) );
  INVX0 U38 ( .INP(n42), .ZN(n2195) );
  INVX0 U39 ( .INP(n54), .ZN(n2170) );
  INVX0 U40 ( .INP(n54), .ZN(n2171) );
  INVX0 U41 ( .INP(n55), .ZN(n2166) );
  INVX0 U42 ( .INP(n55), .ZN(n2167) );
  INVX0 U43 ( .INP(n56), .ZN(n2162) );
  INVX0 U44 ( .INP(n56), .ZN(n2163) );
  INVX0 U45 ( .INP(n63), .ZN(n2138) );
  INVX0 U46 ( .INP(n63), .ZN(n2139) );
  INVX0 U47 ( .INP(n64), .ZN(n2134) );
  INVX0 U48 ( .INP(n64), .ZN(n2135) );
  INVX0 U49 ( .INP(n65), .ZN(n2130) );
  INVX0 U50 ( .INP(n65), .ZN(n2131) );
  INVX0 U51 ( .INP(n72), .ZN(n2106) );
  INVX0 U52 ( .INP(n72), .ZN(n2107) );
  INVX0 U53 ( .INP(n73), .ZN(n2102) );
  INVX0 U54 ( .INP(n73), .ZN(n2103) );
  INVX0 U55 ( .INP(n74), .ZN(n2098) );
  INVX0 U56 ( .INP(n74), .ZN(n2099) );
  INVX0 U57 ( .INP(n52), .ZN(n2174) );
  INVX0 U58 ( .INP(n52), .ZN(n2175) );
  INVX0 U59 ( .INP(n57), .ZN(n2158) );
  INVX0 U60 ( .INP(n57), .ZN(n2159) );
  INVX0 U61 ( .INP(n58), .ZN(n2154) );
  INVX0 U62 ( .INP(n58), .ZN(n2155) );
  INVX0 U63 ( .INP(n59), .ZN(n2150) );
  INVX0 U64 ( .INP(n59), .ZN(n2151) );
  INVX0 U65 ( .INP(n60), .ZN(n2146) );
  INVX0 U66 ( .INP(n60), .ZN(n2147) );
  INVX0 U67 ( .INP(n61), .ZN(n2142) );
  INVX0 U68 ( .INP(n61), .ZN(n2143) );
  INVX0 U69 ( .INP(n66), .ZN(n2126) );
  INVX0 U70 ( .INP(n66), .ZN(n2127) );
  INVX0 U71 ( .INP(n67), .ZN(n2122) );
  INVX0 U72 ( .INP(n67), .ZN(n2123) );
  INVX0 U73 ( .INP(n68), .ZN(n2118) );
  INVX0 U74 ( .INP(n68), .ZN(n2119) );
  INVX0 U75 ( .INP(n69), .ZN(n2114) );
  INVX0 U76 ( .INP(n69), .ZN(n2115) );
  INVX0 U77 ( .INP(n70), .ZN(n2110) );
  INVX0 U78 ( .INP(n70), .ZN(n2111) );
  INVX0 U79 ( .INP(n75), .ZN(n2094) );
  INVX0 U80 ( .INP(n75), .ZN(n2095) );
  INVX0 U81 ( .INP(n76), .ZN(n2090) );
  INVX0 U82 ( .INP(n76), .ZN(n2091) );
  INVX0 U83 ( .INP(n77), .ZN(n2086) );
  INVX0 U84 ( .INP(n77), .ZN(n2087) );
  INVX0 U85 ( .INP(n78), .ZN(n2082) );
  INVX0 U86 ( .INP(n78), .ZN(n2083) );
  INVX0 U87 ( .INP(n44), .ZN(n2190) );
  INVX0 U88 ( .INP(n44), .ZN(n2191) );
  INVX0 U89 ( .INP(n46), .ZN(n2186) );
  INVX0 U90 ( .INP(n46), .ZN(n2187) );
  INVX0 U91 ( .INP(n48), .ZN(n2182) );
  INVX0 U92 ( .INP(n48), .ZN(n2183) );
  INVX0 U93 ( .INP(n50), .ZN(n2178) );
  INVX0 U94 ( .INP(n50), .ZN(n2179) );
  NBUFFX2 U95 ( .INP(n2388), .Z(n2311) );
  NBUFFX2 U96 ( .INP(n2388), .Z(n2312) );
  NBUFFX2 U97 ( .INP(n2388), .Z(n2313) );
  NBUFFX2 U98 ( .INP(n2388), .Z(n2314) );
  NBUFFX2 U99 ( .INP(n2388), .Z(n2315) );
  NBUFFX2 U1104 ( .INP(n2388), .Z(n2316) );
  NBUFFX2 U1105 ( .INP(n2388), .Z(n2317) );
  NBUFFX2 U1106 ( .INP(n2388), .Z(n2318) );
  NBUFFX2 U1107 ( .INP(n2388), .Z(n2319) );
  NBUFFX2 U1108 ( .INP(n2388), .Z(n2320) );
  NBUFFX2 U1109 ( .INP(n2388), .Z(n2321) );
  NBUFFX2 U1110 ( .INP(n2388), .Z(n2322) );
  NBUFFX2 U1111 ( .INP(n2387), .Z(n2323) );
  NBUFFX2 U1112 ( .INP(n2387), .Z(n2324) );
  NBUFFX2 U1113 ( .INP(n2387), .Z(n2325) );
  NBUFFX2 U1114 ( .INP(n2387), .Z(n2326) );
  NBUFFX2 U1115 ( .INP(n2387), .Z(n2327) );
  NBUFFX2 U1116 ( .INP(n2387), .Z(n2328) );
  NBUFFX2 U1117 ( .INP(n2387), .Z(n2329) );
  NBUFFX2 U1118 ( .INP(n2387), .Z(n2330) );
  NBUFFX2 U1119 ( .INP(n2387), .Z(n2331) );
  NBUFFX2 U1120 ( .INP(n2387), .Z(n2332) );
  NBUFFX2 U1121 ( .INP(n2387), .Z(n2333) );
  NBUFFX2 U1122 ( .INP(n2387), .Z(n2334) );
  NBUFFX2 U1123 ( .INP(n2386), .Z(n2335) );
  NBUFFX2 U1124 ( .INP(n2386), .Z(n2336) );
  NBUFFX2 U1125 ( .INP(n2386), .Z(n2337) );
  NBUFFX2 U1126 ( .INP(n2386), .Z(n2338) );
  NBUFFX2 U1127 ( .INP(n2386), .Z(n2339) );
  NBUFFX2 U1128 ( .INP(n2386), .Z(n2340) );
  NBUFFX2 U1129 ( .INP(n2386), .Z(n2341) );
  NBUFFX2 U1130 ( .INP(n2386), .Z(n2342) );
  NBUFFX2 U1131 ( .INP(n2386), .Z(n2343) );
  NBUFFX2 U1132 ( .INP(n2386), .Z(n2344) );
  NBUFFX2 U1133 ( .INP(n2386), .Z(n2345) );
  NBUFFX2 U1134 ( .INP(n2386), .Z(n2346) );
  NBUFFX2 U1135 ( .INP(n2385), .Z(n2347) );
  NBUFFX2 U1136 ( .INP(n2385), .Z(n2348) );
  NBUFFX2 U1137 ( .INP(n2385), .Z(n2349) );
  NBUFFX2 U1138 ( .INP(n2385), .Z(n2350) );
  NBUFFX2 U1139 ( .INP(n2385), .Z(n2351) );
  NBUFFX2 U1140 ( .INP(n2385), .Z(n2352) );
  NBUFFX2 U1141 ( .INP(n2385), .Z(n2353) );
  NBUFFX2 U1142 ( .INP(n2385), .Z(n2354) );
  NBUFFX2 U1143 ( .INP(n2385), .Z(n2355) );
  NBUFFX2 U1144 ( .INP(n2385), .Z(n2356) );
  NBUFFX2 U1145 ( .INP(n2385), .Z(n2357) );
  NBUFFX2 U1146 ( .INP(n2385), .Z(n2358) );
  NBUFFX2 U1147 ( .INP(n2384), .Z(n2359) );
  NBUFFX2 U1148 ( .INP(n2384), .Z(n2360) );
  NBUFFX2 U1149 ( .INP(n2384), .Z(n2361) );
  NBUFFX2 U1150 ( .INP(n2384), .Z(n2362) );
  NBUFFX2 U1151 ( .INP(n2384), .Z(n2363) );
  NBUFFX2 U1152 ( .INP(n2384), .Z(n2364) );
  NBUFFX2 U1153 ( .INP(n2384), .Z(n2365) );
  NBUFFX2 U1154 ( .INP(n2384), .Z(n2366) );
  NBUFFX2 U1155 ( .INP(n2384), .Z(n2367) );
  NBUFFX2 U1156 ( .INP(n2384), .Z(n2368) );
  NBUFFX2 U1157 ( .INP(n2384), .Z(n2369) );
  NBUFFX2 U1158 ( .INP(n2384), .Z(n2370) );
  NBUFFX2 U1159 ( .INP(n2383), .Z(n2371) );
  NBUFFX2 U1160 ( .INP(n2383), .Z(n2372) );
  NBUFFX2 U1161 ( .INP(n2383), .Z(n2373) );
  NBUFFX2 U1162 ( .INP(n2383), .Z(n2374) );
  NBUFFX2 U1163 ( .INP(n2383), .Z(n2375) );
  NBUFFX2 U1164 ( .INP(n2383), .Z(n2376) );
  NBUFFX2 U1165 ( .INP(n2383), .Z(n2377) );
  NBUFFX2 U1166 ( .INP(n2383), .Z(n2378) );
  NBUFFX2 U1167 ( .INP(n2383), .Z(n2379) );
  NBUFFX2 U1168 ( .INP(n2383), .Z(n2380) );
  NBUFFX2 U1169 ( .INP(n2383), .Z(n2381) );
  NBUFFX2 U1170 ( .INP(n2389), .Z(n2300) );
  NBUFFX2 U1171 ( .INP(n2389), .Z(n2301) );
  NBUFFX2 U1172 ( .INP(n2389), .Z(n2302) );
  NBUFFX2 U1173 ( .INP(n2389), .Z(n2303) );
  NBUFFX2 U1174 ( .INP(n2389), .Z(n2304) );
  NBUFFX2 U1175 ( .INP(n2389), .Z(n2305) );
  NBUFFX2 U1176 ( .INP(n2389), .Z(n2306) );
  NBUFFX2 U1177 ( .INP(n2389), .Z(n2307) );
  NBUFFX2 U1178 ( .INP(n2389), .Z(n2308) );
  NBUFFX2 U1179 ( .INP(n2389), .Z(n2309) );
  NBUFFX2 U1180 ( .INP(n2389), .Z(n2310) );
  NBUFFX2 U1181 ( .INP(n2383), .Z(n2382) );
  INVX0 U1182 ( .INP(n2047), .ZN(n2079) );
  INVX0 U1183 ( .INP(n1522), .ZN(n1537) );
  INVX0 U1184 ( .INP(n2044), .ZN(n2059) );
  INVX0 U1185 ( .INP(n1525), .ZN(n1557) );
  INVX0 U1186 ( .INP(n2047), .ZN(n2077) );
  INVX0 U1187 ( .INP(n1525), .ZN(n1555) );
  INVX0 U1188 ( .INP(n1525), .ZN(n1556) );
  INVX0 U1189 ( .INP(n2047), .ZN(n2078) );
  NBUFFX2 U1190 ( .INP(rst_n), .Z(n2388) );
  NBUFFX2 U1191 ( .INP(rst_n), .Z(n2387) );
  NBUFFX2 U1192 ( .INP(rst_n), .Z(n2386) );
  NBUFFX2 U1193 ( .INP(rst_n), .Z(n2385) );
  NBUFFX2 U1194 ( .INP(rst_n), .Z(n2384) );
  NBUFFX2 U1195 ( .INP(rst_n), .Z(n2383) );
  NBUFFX2 U1196 ( .INP(rst_n), .Z(n2389) );
  NBUFFX2 U1197 ( .INP(n1521), .Z(n1523) );
  NBUFFX2 U1198 ( .INP(n2043), .Z(n2046) );
  NBUFFX2 U1199 ( .INP(n2042), .Z(n2040) );
  NBUFFX2 U1200 ( .INP(n2042), .Z(n2030) );
  NBUFFX2 U1201 ( .INP(n2044), .Z(n2047) );
  NBUFFX2 U1202 ( .INP(n1521), .Z(n1524) );
  NBUFFX2 U1203 ( .INP(n1521), .Z(n1522) );
  NBUFFX2 U1204 ( .INP(n2043), .Z(n2044) );
  NBUFFX2 U1205 ( .INP(n1520), .Z(n1518) );
  NBUFFX2 U1206 ( .INP(n2041), .Z(n2021) );
  NBUFFX2 U1207 ( .INP(n1520), .Z(n1508) );
  NBUFFX2 U1208 ( .INP(n1520), .Z(n1509) );
  NBUFFX2 U1209 ( .INP(n2042), .Z(n2031) );
  NBUFFX2 U1210 ( .INP(n2042), .Z(n2029) );
  NBUFFX2 U1211 ( .INP(n2041), .Z(n2022) );
  NBUFFX2 U1212 ( .INP(n1522), .Z(n1525) );
  NBUFFX2 U1213 ( .INP(n1522), .Z(n1526) );
  NBUFFX2 U1214 ( .INP(n2044), .Z(n2048) );
  NBUFFX2 U1215 ( .INP(n2044), .Z(n2049) );
  NBUFFX2 U1216 ( .INP(n2042), .Z(n2039) );
  NBUFFX2 U1217 ( .INP(n1520), .Z(n1516) );
  NBUFFX2 U1218 ( .INP(n2042), .Z(n2038) );
  NBUFFX2 U1219 ( .INP(n1520), .Z(n1510) );
  NBUFFX2 U1220 ( .INP(n2042), .Z(n2032) );
  NBUFFX2 U1221 ( .INP(n2042), .Z(n2033) );
  NBUFFX2 U1222 ( .INP(n1519), .Z(n1499) );
  NBUFFX2 U1223 ( .INP(n1519), .Z(n1502) );
  NBUFFX2 U1224 ( .INP(n2041), .Z(n2024) );
  NBUFFX2 U1225 ( .INP(n1520), .Z(n1507) );
  NBUFFX2 U1226 ( .INP(n1519), .Z(n1500) );
  NBUFFX2 U1227 ( .INP(n1522), .Z(n1527) );
  NBUFFX2 U1228 ( .INP(n2049), .Z(n2050) );
  NBUFFX2 U1229 ( .INP(n1520), .Z(n1517) );
  NBUFFX2 U1230 ( .INP(n1520), .Z(n1511) );
  NBUFFX2 U1231 ( .INP(n2042), .Z(n2034) );
  NBUFFX2 U1232 ( .INP(n1527), .Z(n1528) );
  NBUFFX2 U1233 ( .INP(n2049), .Z(n2051) );
  NBUFFX2 U1234 ( .INP(n1520), .Z(n1512) );
  NBUFFX2 U1235 ( .INP(n1520), .Z(n1513) );
  NBUFFX2 U1236 ( .INP(n2042), .Z(n2035) );
  NBUFFX2 U1237 ( .INP(n2042), .Z(n2036) );
  NBUFFX2 U1238 ( .INP(n1527), .Z(n1529) );
  NBUFFX2 U1239 ( .INP(n2049), .Z(n2052) );
  NBUFFX2 U1240 ( .INP(n1520), .Z(n1514) );
  NBUFFX2 U1241 ( .INP(n1520), .Z(n1515) );
  NBUFFX2 U1242 ( .INP(n2042), .Z(n2037) );
  NBUFFX2 U1243 ( .INP(n2041), .Z(n2023) );
  NBUFFX2 U1244 ( .INP(n1527), .Z(n1530) );
  NBUFFX2 U1245 ( .INP(n1530), .Z(n1531) );
  NBUFFX2 U1246 ( .INP(n2052), .Z(n2053) );
  NBUFFX2 U1247 ( .INP(n2052), .Z(n2054) );
  INVX0 U1248 ( .INP(wr_addr[0]), .ZN(n2390) );
  INVX0 U1249 ( .INP(wr_addr[1]), .ZN(n2391) );
  INVX0 U1250 ( .INP(wr_addr[4]), .ZN(n2393) );
  INVX0 U1251 ( .INP(wr_addr[3]), .ZN(n2392) );
  NBUFFX2 U1252 ( .INP(n2041), .Z(n2025) );
  NBUFFX2 U1253 ( .INP(n2041), .Z(n2026) );
  NBUFFX2 U1254 ( .INP(n1519), .Z(n1501) );
  NBUFFX2 U1255 ( .INP(n1530), .Z(n1532) );
  NBUFFX2 U1256 ( .INP(n2052), .Z(n2055) );
  NBUFFX2 U1257 ( .INP(n1519), .Z(n1503) );
  NBUFFX2 U1258 ( .INP(n1519), .Z(n1504) );
  NBUFFX2 U1259 ( .INP(n2041), .Z(n2027) );
  NBUFFX2 U1260 ( .INP(n1530), .Z(n1533) );
  NBUFFX2 U1261 ( .INP(n2055), .Z(n2056) );
  NBUFFX2 U1262 ( .INP(n1519), .Z(n1505) );
  NBUFFX2 U1263 ( .INP(n2041), .Z(n2028) );
  NBUFFX2 U1264 ( .INP(n1533), .Z(n1534) );
  NBUFFX2 U1265 ( .INP(n2055), .Z(n2057) );
  NBUFFX2 U1266 ( .INP(n1519), .Z(n1506) );
  NBUFFX2 U1267 ( .INP(n1533), .Z(n1535) );
  NAND2X1 U1268 ( .IN1(n2062), .IN2(reg2[1]), .QN(n1998) );
  NAND2X1 U1269 ( .IN1(n1540), .IN2(reg2[1]), .QN(n1476) );
  NAND2X1 U1270 ( .IN1(n2062), .IN2(reg2[2]), .QN(n1994) );
  NAND2X1 U1271 ( .IN1(n2062), .IN2(reg2[3]), .QN(n1990) );
  NAND2X1 U1272 ( .IN1(n2061), .IN2(reg2[4]), .QN(n1986) );
  NAND2X1 U1273 ( .IN1(n1989), .IN2(n1988), .QN(n1606) );
  NAND2X1 U1274 ( .IN1(reg3[4]), .IN2(n2048), .QN(n1987) );
  NAND2X1 U1275 ( .IN1(n2001), .IN2(n2000), .QN(n1576) );
  NAND2X1 U1276 ( .IN1(reg3[1]), .IN2(n2047), .QN(n1999) );
  NAND2X1 U1277 ( .IN1(n1479), .IN2(n1478), .QN(n19) );
  NAND2X1 U1278 ( .IN1(reg3[1]), .IN2(n1525), .QN(n1477) );
  NAND2X1 U1279 ( .IN1(n1997), .IN2(n1996), .QN(n1586) );
  NAND2X1 U1280 ( .IN1(reg3[2]), .IN2(n2048), .QN(n1995) );
  NAND2X1 U1281 ( .IN1(n1993), .IN2(n1992), .QN(n1596) );
  NAND2X1 U1282 ( .IN1(reg3[3]), .IN2(n2048), .QN(n1991) );
  NAND2X1 U1283 ( .IN1(n1540), .IN2(reg2[0]), .QN(n1480) );
  NAND2X1 U1284 ( .IN1(n1540), .IN2(reg2[2]), .QN(n1472) );
  NAND2X1 U1285 ( .IN1(n1540), .IN2(reg2[3]), .QN(n1468) );
  NAND2X1 U1286 ( .IN1(n2062), .IN2(reg2[0]), .QN(n2002) );
  NAND2X1 U1287 ( .IN1(n1539), .IN2(reg2[4]), .QN(n1464) );
  NAND2X1 U1288 ( .IN1(n2061), .IN2(reg2[5]), .QN(n1982) );
  NAND2X1 U1289 ( .IN1(n2061), .IN2(reg2[6]), .QN(n1978) );
  NAND2X1 U1290 ( .IN1(n2061), .IN2(reg2[7]), .QN(n1974) );
  NAND2X1 U1291 ( .IN1(n1467), .IN2(n1466), .QN(n1084) );
  NAND2X1 U1292 ( .IN1(reg3[4]), .IN2(n1526), .QN(n1465) );
  NAND2X1 U1293 ( .IN1(n1985), .IN2(n1984), .QN(n1616) );
  NAND2X1 U1294 ( .IN1(reg3[5]), .IN2(n2049), .QN(n1983) );
  NAND2X1 U1295 ( .IN1(n1981), .IN2(n1980), .QN(n1626) );
  NAND2X1 U1296 ( .IN1(reg3[6]), .IN2(n2049), .QN(n1979) );
  NAND2X1 U1297 ( .IN1(n1977), .IN2(n1976), .QN(n1636) );
  NAND2X1 U1298 ( .IN1(reg3[7]), .IN2(n2049), .QN(n1975) );
  NAND2X1 U1299 ( .IN1(n1483), .IN2(n1482), .QN(n9) );
  NAND2X1 U1300 ( .IN1(reg3[0]), .IN2(n1525), .QN(n1481) );
  NAND2X1 U1301 ( .IN1(n2005), .IN2(n2004), .QN(n1566) );
  NAND2X1 U1302 ( .IN1(reg3[0]), .IN2(n2047), .QN(n2003) );
  NAND2X1 U1303 ( .IN1(n1475), .IN2(n1474), .QN(n29) );
  NAND2X1 U1304 ( .IN1(reg3[2]), .IN2(n1526), .QN(n1473) );
  NAND2X1 U1305 ( .IN1(n1471), .IN2(n1470), .QN(n1074) );
  NAND2X1 U1306 ( .IN1(reg3[3]), .IN2(n1526), .QN(n1469) );
  NAND2X1 U1307 ( .IN1(n1539), .IN2(reg2[5]), .QN(n1460) );
  NAND2X1 U1308 ( .IN1(n1539), .IN2(reg2[6]), .QN(n1456) );
  NAND2X1 U1309 ( .IN1(n1539), .IN2(reg2[7]), .QN(n1452) );
  NAND2X1 U1310 ( .IN1(n1539), .IN2(reg2[8]), .QN(n1448) );
  NAND2X1 U1311 ( .IN1(n2061), .IN2(reg2[8]), .QN(n1970) );
  NAND2X1 U1312 ( .IN1(n2061), .IN2(reg2[9]), .QN(n1966) );
  NAND2X1 U1313 ( .IN1(n2061), .IN2(reg2[10]), .QN(n1962) );
  NAND2X1 U1314 ( .IN1(n2061), .IN2(reg2[11]), .QN(n1958) );
  NBUFFX2 U1315 ( .INP(N17), .Z(n2042) );
  NAND2X1 U1316 ( .IN1(n1463), .IN2(n1462), .QN(n1094) );
  NAND2X1 U1317 ( .IN1(reg3[5]), .IN2(n1527), .QN(n1461) );
  NAND2X1 U1318 ( .IN1(n1459), .IN2(n1458), .QN(n1104) );
  NAND2X1 U1319 ( .IN1(reg3[6]), .IN2(n1527), .QN(n1457) );
  NAND2X1 U1320 ( .IN1(n1455), .IN2(n1454), .QN(n1114) );
  NAND2X1 U1321 ( .IN1(reg3[7]), .IN2(n1527), .QN(n1453) );
  NAND2X1 U1322 ( .IN1(n1451), .IN2(n1450), .QN(n1124) );
  NAND2X1 U1323 ( .IN1(reg3[8]), .IN2(n1528), .QN(n1449) );
  NAND2X1 U1324 ( .IN1(n1973), .IN2(n1972), .QN(n1646) );
  NAND2X1 U1325 ( .IN1(reg3[8]), .IN2(n2050), .QN(n1971) );
  NAND2X1 U1326 ( .IN1(n1969), .IN2(n1968), .QN(n1656) );
  NAND2X1 U1327 ( .IN1(reg3[9]), .IN2(n2050), .QN(n1967) );
  NAND2X1 U1328 ( .IN1(n1965), .IN2(n1964), .QN(n1666) );
  NAND2X1 U1329 ( .IN1(reg3[10]), .IN2(n2050), .QN(n1963) );
  NAND2X1 U1330 ( .IN1(n1961), .IN2(n1960), .QN(n1676) );
  NAND2X1 U1331 ( .IN1(reg3[11]), .IN2(n2051), .QN(n1959) );
  NAND2X1 U1332 ( .IN1(n1539), .IN2(reg2[9]), .QN(n1444) );
  NAND2X1 U1333 ( .IN1(n1539), .IN2(reg2[10]), .QN(n1440) );
  NAND2X1 U1334 ( .IN1(n1539), .IN2(reg2[11]), .QN(n1436) );
  NAND2X1 U1335 ( .IN1(n1539), .IN2(reg2[12]), .QN(n1432) );
  NAND2X1 U1336 ( .IN1(n2061), .IN2(reg2[12]), .QN(n1954) );
  NAND2X1 U1337 ( .IN1(n2061), .IN2(reg2[13]), .QN(n1950) );
  NAND2X1 U1338 ( .IN1(n2061), .IN2(reg2[14]), .QN(n1946) );
  NAND2X1 U1339 ( .IN1(n2061), .IN2(reg2[15]), .QN(n1942) );
  NBUFFX2 U1340 ( .INP(N17), .Z(n2041) );
  NBUFFX2 U1341 ( .INP(N12), .Z(n1520) );
  NAND2X1 U1342 ( .IN1(n1447), .IN2(n1446), .QN(n1134) );
  NAND2X1 U1343 ( .IN1(reg3[9]), .IN2(n1528), .QN(n1445) );
  NAND2X1 U1344 ( .IN1(n1443), .IN2(n1442), .QN(n1144) );
  NAND2X1 U1345 ( .IN1(reg3[10]), .IN2(n1528), .QN(n1441) );
  NAND2X1 U1346 ( .IN1(n1439), .IN2(n1438), .QN(n1154) );
  NAND2X1 U1347 ( .IN1(reg3[11]), .IN2(n1529), .QN(n1437) );
  NAND2X1 U1348 ( .IN1(n1435), .IN2(n1434), .QN(n1164) );
  NAND2X1 U1349 ( .IN1(reg3[12]), .IN2(n1529), .QN(n1433) );
  NAND2X1 U1350 ( .IN1(n1957), .IN2(n1956), .QN(n1686) );
  NAND2X1 U1351 ( .IN1(reg3[12]), .IN2(n2051), .QN(n1955) );
  NAND2X1 U1352 ( .IN1(n1953), .IN2(n1952), .QN(n1696) );
  NAND2X1 U1353 ( .IN1(reg3[13]), .IN2(n2051), .QN(n1951) );
  NAND2X1 U1354 ( .IN1(n1949), .IN2(n1948), .QN(n1706) );
  NAND2X1 U1355 ( .IN1(reg3[14]), .IN2(n2052), .QN(n1947) );
  NAND2X1 U1356 ( .IN1(n1945), .IN2(n1944), .QN(n1716) );
  NAND2X1 U1357 ( .IN1(reg3[15]), .IN2(n2052), .QN(n1943) );
  NBUFFX4 U1358 ( .INP(N13), .Z(n1494) );
  NBUFFX4 U1359 ( .INP(N18), .Z(n2016) );
  NAND2X1 U1360 ( .IN1(n1539), .IN2(reg2[13]), .QN(n1428) );
  NAND2X1 U1361 ( .IN1(n1539), .IN2(reg2[14]), .QN(n1424) );
  NAND2X1 U1362 ( .IN1(n1539), .IN2(reg2[15]), .QN(n1420) );
  NAND2X1 U1363 ( .IN1(n1539), .IN2(reg2[16]), .QN(n1416) );
  NAND2X1 U1364 ( .IN1(n2061), .IN2(reg2[16]), .QN(n1938) );
  NAND2X1 U1365 ( .IN1(n2060), .IN2(reg2[17]), .QN(n1934) );
  NAND2X1 U1366 ( .IN1(n2060), .IN2(reg2[18]), .QN(n1930) );
  NAND2X1 U1367 ( .IN1(n2060), .IN2(reg2[19]), .QN(n1926) );
  NBUFFX2 U1368 ( .INP(N12), .Z(n1519) );
  NAND2X1 U1369 ( .IN1(n1431), .IN2(n1430), .QN(n1174) );
  NAND2X1 U1370 ( .IN1(reg3[13]), .IN2(n1529), .QN(n1429) );
  NAND2X1 U1371 ( .IN1(n1427), .IN2(n1426), .QN(n1184) );
  NAND2X1 U1372 ( .IN1(reg3[14]), .IN2(n1530), .QN(n1425) );
  NAND2X1 U1373 ( .IN1(n1423), .IN2(n1422), .QN(n1194) );
  NAND2X1 U1374 ( .IN1(reg3[15]), .IN2(n1530), .QN(n1421) );
  NAND2X1 U1375 ( .IN1(n1419), .IN2(n1418), .QN(n1204) );
  NAND2X1 U1376 ( .IN1(reg3[16]), .IN2(n1530), .QN(n1417) );
  NAND2X1 U1377 ( .IN1(n1941), .IN2(n1940), .QN(n1726) );
  NAND2X1 U1378 ( .IN1(reg3[16]), .IN2(n2052), .QN(n1939) );
  NAND2X1 U1379 ( .IN1(n1937), .IN2(n1936), .QN(n1736) );
  NAND2X1 U1380 ( .IN1(reg3[17]), .IN2(n2053), .QN(n1935) );
  NAND2X1 U1381 ( .IN1(n1933), .IN2(n1932), .QN(n1746) );
  NAND2X1 U1382 ( .IN1(reg3[18]), .IN2(n2053), .QN(n1931) );
  NAND2X1 U1383 ( .IN1(n1929), .IN2(n1928), .QN(n1756) );
  NAND2X1 U1384 ( .IN1(reg3[19]), .IN2(n2053), .QN(n1927) );
  NBUFFX4 U1385 ( .INP(N18), .Z(n2017) );
  NBUFFX2 U1386 ( .INP(N19), .Z(n2009) );
  NAND2X1 U1387 ( .IN1(n1538), .IN2(reg2[17]), .QN(n1412) );
  NAND2X1 U1388 ( .IN1(n1538), .IN2(reg2[18]), .QN(n1408) );
  NAND2X1 U1389 ( .IN1(n1538), .IN2(reg2[19]), .QN(n1404) );
  NAND2X1 U1390 ( .IN1(n2060), .IN2(reg2[20]), .QN(n1922) );
  NAND2X1 U1391 ( .IN1(n2060), .IN2(reg2[21]), .QN(n1918) );
  NAND2X1 U1392 ( .IN1(n2060), .IN2(reg2[22]), .QN(n1914) );
  NBUFFX2 U1393 ( .INP(N19), .Z(n2010) );
  NBUFFX2 U1394 ( .INP(N20), .Z(n2006) );
  NBUFFX2 U1395 ( .INP(N13), .Z(n1493) );
  NBUFFX2 U1396 ( .INP(N18), .Z(n2015) );
  NAND2X1 U1397 ( .IN1(n2059), .IN2(reg2[30]), .QN(n1882) );
  NAND2X1 U1398 ( .IN1(n1415), .IN2(n1414), .QN(n1214) );
  NAND2X1 U1399 ( .IN1(reg3[17]), .IN2(n1531), .QN(n1413) );
  NAND2X1 U1400 ( .IN1(n1411), .IN2(n1410), .QN(n1224) );
  NAND2X1 U1401 ( .IN1(reg3[18]), .IN2(n1531), .QN(n1409) );
  NAND2X1 U1402 ( .IN1(n1407), .IN2(n1406), .QN(n1234) );
  NAND2X1 U1403 ( .IN1(reg3[19]), .IN2(n1531), .QN(n1405) );
  NAND2X1 U1404 ( .IN1(n1925), .IN2(n1924), .QN(n1766) );
  NAND2X1 U1405 ( .IN1(reg3[20]), .IN2(n2054), .QN(n1923) );
  NAND2X1 U1406 ( .IN1(n1921), .IN2(n1920), .QN(n1776) );
  NAND2X1 U1407 ( .IN1(reg3[21]), .IN2(n2054), .QN(n1919) );
  NAND2X1 U1408 ( .IN1(n1917), .IN2(n1916), .QN(n1786) );
  NAND2X1 U1409 ( .IN1(reg3[22]), .IN2(n2054), .QN(n1915) );
  NAND2X1 U1410 ( .IN1(n1885), .IN2(n1884), .QN(n1866) );
  NAND2X1 U1411 ( .IN1(reg3[30]), .IN2(n2057), .QN(n1883) );
  NBUFFX4 U1412 ( .INP(N13), .Z(n1495) );
  NBUFFX2 U1413 ( .INP(N14), .Z(n1487) );
  NAND2X1 U1414 ( .IN1(n1538), .IN2(reg2[20]), .QN(n1400) );
  NAND2X1 U1415 ( .IN1(n1538), .IN2(reg2[21]), .QN(n1396) );
  NAND2X1 U1416 ( .IN1(n1538), .IN2(reg2[22]), .QN(n1392) );
  NAND2X1 U1417 ( .IN1(n1538), .IN2(reg2[23]), .QN(n1388) );
  NAND2X1 U1418 ( .IN1(n2060), .IN2(reg2[23]), .QN(n1910) );
  NAND2X1 U1419 ( .IN1(n2060), .IN2(reg2[24]), .QN(n1906) );
  NAND2X1 U1420 ( .IN1(n2060), .IN2(reg2[25]), .QN(n1902) );
  NAND2X1 U1421 ( .IN1(n2060), .IN2(reg2[26]), .QN(n1898) );
  NBUFFX2 U1422 ( .INP(N14), .Z(n1488) );
  NBUFFX2 U1423 ( .INP(N19), .Z(n2011) );
  NBUFFX2 U1424 ( .INP(N15), .Z(n1484) );
  NAND2X1 U1425 ( .IN1(n1537), .IN2(reg2[30]), .QN(n1360) );
  NAND2X1 U1426 ( .IN1(n1403), .IN2(n1402), .QN(n1244) );
  NAND2X1 U1427 ( .IN1(reg3[20]), .IN2(n1532), .QN(n1401) );
  NAND2X1 U1428 ( .IN1(n1399), .IN2(n1398), .QN(n1254) );
  NAND2X1 U1429 ( .IN1(reg3[21]), .IN2(n1532), .QN(n1397) );
  NAND2X1 U1430 ( .IN1(n1395), .IN2(n1394), .QN(n1264) );
  NAND2X1 U1431 ( .IN1(reg3[22]), .IN2(n1532), .QN(n1393) );
  NAND2X1 U1432 ( .IN1(n1391), .IN2(n1390), .QN(n1274) );
  NAND2X1 U1433 ( .IN1(reg3[23]), .IN2(n1533), .QN(n1389) );
  NAND2X1 U1434 ( .IN1(n1913), .IN2(n1912), .QN(n1796) );
  NAND2X1 U1435 ( .IN1(reg3[23]), .IN2(n2055), .QN(n1911) );
  NAND2X1 U1436 ( .IN1(n1909), .IN2(n1908), .QN(n1806) );
  NAND2X1 U1437 ( .IN1(reg3[24]), .IN2(n2055), .QN(n1907) );
  NAND2X1 U1438 ( .IN1(n1905), .IN2(n1904), .QN(n1816) );
  NAND2X1 U1439 ( .IN1(reg3[25]), .IN2(n2055), .QN(n1903) );
  NAND2X1 U1440 ( .IN1(n1901), .IN2(n1900), .QN(n1826) );
  NAND2X1 U1441 ( .IN1(reg3[26]), .IN2(n2056), .QN(n1899) );
  NAND2X1 U1442 ( .IN1(n1363), .IN2(n1362), .QN(n1344) );
  NAND2X1 U1443 ( .IN1(reg3[30]), .IN2(n1535), .QN(n1361) );
  NBUFFX4 U1444 ( .INP(N18), .Z(n2018) );
  NBUFFX2 U1445 ( .INP(N20), .Z(n2007) );
  NAND2X1 U1446 ( .IN1(n1538), .IN2(reg2[24]), .QN(n1384) );
  NAND2X1 U1447 ( .IN1(n1538), .IN2(reg2[25]), .QN(n1380) );
  NAND2X1 U1448 ( .IN1(n1538), .IN2(reg2[26]), .QN(n1376) );
  NAND2X1 U1449 ( .IN1(n1538), .IN2(reg2[27]), .QN(n1372) );
  NAND2X1 U1450 ( .IN1(n2060), .IN2(reg2[27]), .QN(n1894) );
  NAND2X1 U1451 ( .IN1(n2060), .IN2(reg2[28]), .QN(n1890) );
  NAND2X1 U1452 ( .IN1(n2060), .IN2(reg2[29]), .QN(n1886) );
  NBUFFX2 U1453 ( .INP(N14), .Z(n1489) );
  NAND2X1 U1454 ( .IN1(n1387), .IN2(n1386), .QN(n1284) );
  NAND2X1 U1455 ( .IN1(reg3[24]), .IN2(n1533), .QN(n1385) );
  NAND2X1 U1456 ( .IN1(n1383), .IN2(n1382), .QN(n1294) );
  NAND2X1 U1457 ( .IN1(reg3[25]), .IN2(n1533), .QN(n1381) );
  NAND2X1 U1458 ( .IN1(n1379), .IN2(n1378), .QN(n1304) );
  NAND2X1 U1459 ( .IN1(reg3[26]), .IN2(n1534), .QN(n1377) );
  NAND2X1 U1460 ( .IN1(n1375), .IN2(n1374), .QN(n1314) );
  NAND2X1 U1461 ( .IN1(reg3[27]), .IN2(n1534), .QN(n1373) );
  NAND2X1 U1462 ( .IN1(n1897), .IN2(n1896), .QN(n1836) );
  NAND2X1 U1463 ( .IN1(reg3[27]), .IN2(n2056), .QN(n1895) );
  NAND2X1 U1464 ( .IN1(n1893), .IN2(n1892), .QN(n1846) );
  NAND2X1 U1465 ( .IN1(reg3[28]), .IN2(n2056), .QN(n1891) );
  NAND2X1 U1466 ( .IN1(n1889), .IN2(n1888), .QN(n1856) );
  NAND2X1 U1467 ( .IN1(reg3[29]), .IN2(n2057), .QN(n1887) );
  NBUFFX4 U1468 ( .INP(N13), .Z(n1496) );
  NBUFFX4 U1469 ( .INP(N18), .Z(n2019) );
  NAND2X1 U1470 ( .IN1(n2062), .IN2(reg2[31]), .QN(n1878) );
  NBUFFX2 U1471 ( .INP(N15), .Z(n1485) );
  NAND2X1 U1472 ( .IN1(n1538), .IN2(reg2[28]), .QN(n1368) );
  NAND2X1 U1473 ( .IN1(n1538), .IN2(reg2[29]), .QN(n1364) );
  NBUFFX2 U1474 ( .INP(N19), .Z(n2012) );
  NAND2X1 U1475 ( .IN1(n1371), .IN2(n1370), .QN(n1324) );
  NAND2X1 U1476 ( .IN1(reg3[28]), .IN2(n1534), .QN(n1369) );
  NAND2X1 U1477 ( .IN1(n1367), .IN2(n1366), .QN(n1334) );
  NAND2X1 U1478 ( .IN1(reg3[29]), .IN2(n1535), .QN(n1365) );
  NAND2X1 U1479 ( .IN1(n1881), .IN2(n1880), .QN(n1876) );
  NAND2X1 U1480 ( .IN1(reg3[31]), .IN2(n2057), .QN(n1879) );
  NBUFFX4 U1481 ( .INP(N13), .Z(n1497) );
  NAND2X1 U1482 ( .IN1(n1540), .IN2(reg2[31]), .QN(n1356) );
  NBUFFX2 U1483 ( .INP(N14), .Z(n1490) );
  NAND2X1 U1484 ( .IN1(n1359), .IN2(n1358), .QN(n1354) );
  NAND2X1 U1485 ( .IN1(reg3[31]), .IN2(n1535), .QN(n1357) );
  NBUFFX4 U1486 ( .INP(N18), .Z(n2020) );
  NBUFFX2 U1487 ( .INP(N20), .Z(n2008) );
  NBUFFX2 U1488 ( .INP(N14), .Z(n1491) );
  NBUFFX2 U1489 ( .INP(N19), .Z(n2013) );
  NBUFFX4 U1490 ( .INP(N13), .Z(n1498) );
  NBUFFX2 U1491 ( .INP(N15), .Z(n1486) );
  NBUFFX2 U1492 ( .INP(N19), .Z(n2014) );
  NBUFFX2 U1493 ( .INP(N14), .Z(n1492) );
  NBUFFX2 U1494 ( .INP(wr_data[0]), .Z(n2204) );
  NBUFFX2 U1495 ( .INP(wr_data[1]), .Z(n2207) );
  NBUFFX2 U1496 ( .INP(wr_data[2]), .Z(n2210) );
  NBUFFX2 U1497 ( .INP(wr_data[3]), .Z(n2213) );
  NBUFFX2 U1498 ( .INP(wr_data[4]), .Z(n2216) );
  NBUFFX2 U1499 ( .INP(wr_data[5]), .Z(n2219) );
  NBUFFX2 U1500 ( .INP(wr_data[6]), .Z(n2222) );
  NBUFFX2 U1501 ( .INP(wr_data[7]), .Z(n2225) );
  NBUFFX2 U1502 ( .INP(wr_data[8]), .Z(n2228) );
  NBUFFX2 U1503 ( .INP(wr_data[9]), .Z(n2231) );
  NBUFFX2 U1504 ( .INP(wr_data[10]), .Z(n2234) );
  NBUFFX2 U1505 ( .INP(wr_data[11]), .Z(n2237) );
  NBUFFX2 U1506 ( .INP(wr_data[12]), .Z(n2240) );
  NBUFFX2 U1507 ( .INP(wr_data[13]), .Z(n2243) );
  NBUFFX2 U1508 ( .INP(wr_data[14]), .Z(n2246) );
  NBUFFX2 U1509 ( .INP(wr_data[15]), .Z(n2249) );
  NBUFFX2 U1510 ( .INP(wr_data[16]), .Z(n2252) );
  NBUFFX2 U1511 ( .INP(wr_data[17]), .Z(n2255) );
  NBUFFX2 U1512 ( .INP(wr_data[18]), .Z(n2258) );
  NBUFFX2 U1513 ( .INP(wr_data[19]), .Z(n2261) );
  NBUFFX2 U1514 ( .INP(wr_data[20]), .Z(n2264) );
  NBUFFX2 U1515 ( .INP(wr_data[21]), .Z(n2267) );
  NBUFFX2 U1516 ( .INP(wr_data[22]), .Z(n2270) );
  NBUFFX2 U1517 ( .INP(wr_data[23]), .Z(n2273) );
  NBUFFX2 U1518 ( .INP(wr_data[24]), .Z(n2276) );
  NBUFFX2 U1519 ( .INP(wr_data[25]), .Z(n2279) );
  NBUFFX2 U1520 ( .INP(wr_data[26]), .Z(n2282) );
  NBUFFX2 U1521 ( .INP(wr_data[27]), .Z(n2285) );
  NBUFFX2 U1522 ( .INP(wr_data[28]), .Z(n2288) );
  NBUFFX2 U1523 ( .INP(wr_data[29]), .Z(n2291) );
  NBUFFX2 U1524 ( .INP(wr_data[30]), .Z(n2294) );
  NBUFFX2 U1525 ( .INP(wr_data[31]), .Z(n2297) );
  NBUFFX2 U1526 ( .INP(wr_data[0]), .Z(n2205) );
  NBUFFX2 U1527 ( .INP(wr_data[1]), .Z(n2208) );
  NBUFFX2 U1528 ( .INP(wr_data[2]), .Z(n2211) );
  NBUFFX2 U1529 ( .INP(wr_data[3]), .Z(n2214) );
  NBUFFX2 U1530 ( .INP(wr_data[4]), .Z(n2217) );
  NBUFFX2 U1531 ( .INP(wr_data[5]), .Z(n2220) );
  NBUFFX2 U1532 ( .INP(wr_data[6]), .Z(n2223) );
  NBUFFX2 U1533 ( .INP(wr_data[7]), .Z(n2226) );
  NBUFFX2 U1534 ( .INP(wr_data[8]), .Z(n2229) );
  NBUFFX2 U1535 ( .INP(wr_data[9]), .Z(n2232) );
  NBUFFX2 U1536 ( .INP(wr_data[10]), .Z(n2235) );
  NBUFFX2 U1537 ( .INP(wr_data[11]), .Z(n2238) );
  NBUFFX2 U1538 ( .INP(wr_data[12]), .Z(n2241) );
  NBUFFX2 U1539 ( .INP(wr_data[13]), .Z(n2244) );
  NBUFFX2 U1540 ( .INP(wr_data[14]), .Z(n2247) );
  NBUFFX2 U1541 ( .INP(wr_data[15]), .Z(n2250) );
  NBUFFX2 U1542 ( .INP(wr_data[16]), .Z(n2253) );
  NBUFFX2 U1543 ( .INP(wr_data[17]), .Z(n2256) );
  NBUFFX2 U1544 ( .INP(wr_data[18]), .Z(n2259) );
  NBUFFX2 U1545 ( .INP(wr_data[19]), .Z(n2262) );
  NBUFFX2 U1546 ( .INP(wr_data[20]), .Z(n2265) );
  NBUFFX2 U1547 ( .INP(wr_data[21]), .Z(n2268) );
  NBUFFX2 U1548 ( .INP(wr_data[22]), .Z(n2271) );
  NBUFFX2 U1549 ( .INP(wr_data[23]), .Z(n2274) );
  NBUFFX2 U1550 ( .INP(wr_data[24]), .Z(n2277) );
  NBUFFX2 U1551 ( .INP(wr_data[25]), .Z(n2280) );
  NBUFFX2 U1552 ( .INP(wr_data[26]), .Z(n2283) );
  NBUFFX2 U1553 ( .INP(wr_data[27]), .Z(n2286) );
  NBUFFX2 U1554 ( .INP(wr_data[28]), .Z(n2289) );
  NBUFFX2 U1555 ( .INP(wr_data[29]), .Z(n2292) );
  NBUFFX2 U1556 ( .INP(wr_data[30]), .Z(n2295) );
  NBUFFX2 U1557 ( .INP(wr_data[31]), .Z(n2298) );
  NBUFFX2 U1558 ( .INP(wr_data[0]), .Z(n2206) );
  NBUFFX2 U1559 ( .INP(wr_data[1]), .Z(n2209) );
  NBUFFX2 U1560 ( .INP(wr_data[2]), .Z(n2212) );
  NBUFFX2 U1561 ( .INP(wr_data[3]), .Z(n2215) );
  NBUFFX2 U1562 ( .INP(wr_data[4]), .Z(n2218) );
  NBUFFX2 U1563 ( .INP(wr_data[5]), .Z(n2221) );
  NBUFFX2 U1564 ( .INP(wr_data[6]), .Z(n2224) );
  NBUFFX2 U1565 ( .INP(wr_data[7]), .Z(n2227) );
  NBUFFX2 U1566 ( .INP(wr_data[8]), .Z(n2230) );
  NBUFFX2 U1567 ( .INP(wr_data[9]), .Z(n2233) );
  NBUFFX2 U1568 ( .INP(wr_data[10]), .Z(n2236) );
  NBUFFX2 U1569 ( .INP(wr_data[11]), .Z(n2239) );
  NBUFFX2 U1570 ( .INP(wr_data[12]), .Z(n2242) );
  NBUFFX2 U1571 ( .INP(wr_data[13]), .Z(n2245) );
  NBUFFX2 U1572 ( .INP(wr_data[14]), .Z(n2248) );
  NBUFFX2 U1573 ( .INP(wr_data[15]), .Z(n2251) );
  NBUFFX2 U1574 ( .INP(wr_data[16]), .Z(n2254) );
  NBUFFX2 U1575 ( .INP(wr_data[17]), .Z(n2257) );
  NBUFFX2 U1576 ( .INP(wr_data[18]), .Z(n2260) );
  NBUFFX2 U1577 ( .INP(wr_data[19]), .Z(n2263) );
  NBUFFX2 U1578 ( .INP(wr_data[20]), .Z(n2266) );
  NBUFFX2 U1579 ( .INP(wr_data[21]), .Z(n2269) );
  NBUFFX2 U1580 ( .INP(wr_data[22]), .Z(n2272) );
  NBUFFX2 U1581 ( .INP(wr_data[23]), .Z(n2275) );
  NBUFFX2 U1582 ( .INP(wr_data[24]), .Z(n2278) );
  NBUFFX2 U1583 ( .INP(wr_data[25]), .Z(n2281) );
  NBUFFX2 U1584 ( .INP(wr_data[26]), .Z(n2284) );
  NBUFFX2 U1585 ( .INP(wr_data[27]), .Z(n2287) );
  NBUFFX2 U1586 ( .INP(wr_data[28]), .Z(n2290) );
  NBUFFX2 U1587 ( .INP(wr_data[29]), .Z(n2293) );
  NBUFFX2 U1588 ( .INP(wr_data[30]), .Z(n2296) );
  NBUFFX2 U1589 ( .INP(wr_data[31]), .Z(n2299) );
  MUX41X1 U1590 ( .IN1(reg29[0]), .IN3(reg31[0]), .IN2(reg30[0]), .IN4(
        reg32[0]), .S0(n1502), .S1(n1540), .Q(n1) );
  MUX41X1 U1591 ( .IN1(reg25[0]), .IN3(reg27[0]), .IN2(reg26[0]), .IN4(
        reg28[0]), .S0(n1516), .S1(n1557), .Q(n2) );
  MUX41X1 U1592 ( .IN1(reg21[0]), .IN3(reg23[0]), .IN2(reg22[0]), .IN4(
        reg24[0]), .S0(n1507), .S1(n1547), .Q(n3) );
  MUX41X1 U1593 ( .IN1(reg17[0]), .IN3(reg19[0]), .IN2(reg18[0]), .IN4(
        reg20[0]), .S0(n1507), .S1(n1547), .Q(n4) );
  MUX41X1 U1594 ( .IN1(n4), .IN3(n2), .IN2(n3), .IN4(n1), .S0(n1487), .S1(
        n1493), .Q(n5) );
  MUX41X1 U1595 ( .IN1(reg13[0]), .IN3(reg15[0]), .IN2(reg14[0]), .IN4(
        reg16[0]), .S0(n1508), .S1(n1547), .Q(n6) );
  MUX41X1 U1596 ( .IN1(reg9[0]), .IN3(reg11[0]), .IN2(reg10[0]), .IN4(reg12[0]), .S0(n1508), .S1(n1547), .Q(n7) );
  MUX41X1 U1597 ( .IN1(reg5[0]), .IN3(reg7[0]), .IN2(reg6[0]), .IN4(reg8[0]), 
        .S0(n1508), .S1(n1547), .Q(n8) );
  MUX41X1 U1598 ( .IN1(n9), .IN3(n7), .IN2(n8), .IN4(n6), .S0(n1487), .S1(
        n1493), .Q(n10) );
  MUX21X1 U1599 ( .IN1(n10), .IN2(n5), .S(n1484), .Q(rd_dataA[0]) );
  MUX41X1 U1600 ( .IN1(reg29[1]), .IN3(reg31[1]), .IN2(reg30[1]), .IN4(
        reg32[1]), .S0(n1508), .S1(n1547), .Q(n11) );
  MUX41X1 U1601 ( .IN1(reg25[1]), .IN3(reg27[1]), .IN2(reg26[1]), .IN4(
        reg28[1]), .S0(n1508), .S1(n1547), .Q(n12) );
  MUX41X1 U1602 ( .IN1(reg21[1]), .IN3(reg23[1]), .IN2(reg22[1]), .IN4(
        reg24[1]), .S0(n1508), .S1(n1547), .Q(n13) );
  MUX41X1 U1603 ( .IN1(reg17[1]), .IN3(reg19[1]), .IN2(reg18[1]), .IN4(
        reg20[1]), .S0(n1508), .S1(n1547), .Q(n14) );
  MUX41X1 U1604 ( .IN1(n14), .IN3(n12), .IN2(n13), .IN4(n11), .S0(n1487), .S1(
        n1493), .Q(n15) );
  MUX41X1 U1605 ( .IN1(reg13[1]), .IN3(reg15[1]), .IN2(reg14[1]), .IN4(
        reg16[1]), .S0(n1508), .S1(n1547), .Q(n16) );
  MUX41X1 U1606 ( .IN1(reg9[1]), .IN3(reg11[1]), .IN2(reg10[1]), .IN4(reg12[1]), .S0(n1508), .S1(n1547), .Q(n17) );
  MUX41X1 U1607 ( .IN1(reg5[1]), .IN3(reg7[1]), .IN2(reg6[1]), .IN4(reg8[1]), 
        .S0(n1508), .S1(n1548), .Q(n18) );
  MUX41X1 U1608 ( .IN1(n19), .IN3(n17), .IN2(n18), .IN4(n16), .S0(n1487), .S1(
        n1493), .Q(n20) );
  MUX21X1 U1609 ( .IN1(n20), .IN2(n15), .S(n1484), .Q(rd_dataA[1]) );
  MUX41X1 U1610 ( .IN1(reg29[2]), .IN3(reg31[2]), .IN2(reg30[2]), .IN4(
        reg32[2]), .S0(n1508), .S1(n1548), .Q(n21) );
  MUX41X1 U1611 ( .IN1(reg25[2]), .IN3(reg27[2]), .IN2(reg26[2]), .IN4(
        reg28[2]), .S0(n1508), .S1(n1548), .Q(n22) );
  MUX41X1 U1612 ( .IN1(reg21[2]), .IN3(reg23[2]), .IN2(reg22[2]), .IN4(
        reg24[2]), .S0(n1508), .S1(n1548), .Q(n23) );
  MUX41X1 U1613 ( .IN1(reg17[2]), .IN3(reg19[2]), .IN2(reg18[2]), .IN4(
        reg20[2]), .S0(n1508), .S1(n1548), .Q(n24) );
  MUX41X1 U1614 ( .IN1(n24), .IN3(n22), .IN2(n23), .IN4(n21), .S0(n1488), .S1(
        n1494), .Q(n25) );
  MUX41X1 U1615 ( .IN1(reg13[2]), .IN3(reg15[2]), .IN2(reg14[2]), .IN4(
        reg16[2]), .S0(n1508), .S1(n1548), .Q(n26) );
  MUX41X1 U1616 ( .IN1(reg9[2]), .IN3(reg11[2]), .IN2(reg10[2]), .IN4(reg12[2]), .S0(n1509), .S1(n1548), .Q(n27) );
  MUX41X1 U1617 ( .IN1(reg5[2]), .IN3(reg7[2]), .IN2(reg6[2]), .IN4(reg8[2]), 
        .S0(n1509), .S1(n1548), .Q(n28) );
  MUX41X1 U1618 ( .IN1(n29), .IN3(n27), .IN2(n28), .IN4(n26), .S0(n1488), .S1(
        n1494), .Q(n30) );
  MUX21X1 U1619 ( .IN1(n30), .IN2(n25), .S(n1484), .Q(rd_dataA[2]) );
  MUX41X1 U1620 ( .IN1(reg29[3]), .IN3(reg31[3]), .IN2(reg30[3]), .IN4(
        reg32[3]), .S0(n1509), .S1(n1548), .Q(n31) );
  MUX41X1 U1621 ( .IN1(reg25[3]), .IN3(reg27[3]), .IN2(reg26[3]), .IN4(
        reg28[3]), .S0(n1509), .S1(n1548), .Q(n32) );
  MUX41X1 U1622 ( .IN1(reg21[3]), .IN3(reg23[3]), .IN2(reg22[3]), .IN4(
        reg24[3]), .S0(n1509), .S1(n1548), .Q(n33) );
  MUX41X1 U1623 ( .IN1(reg17[3]), .IN3(reg19[3]), .IN2(reg18[3]), .IN4(
        reg20[3]), .S0(n1509), .S1(n1548), .Q(n34) );
  MUX41X1 U1624 ( .IN1(n34), .IN3(n32), .IN2(n33), .IN4(n31), .S0(n1488), .S1(
        n1494), .Q(n35) );
  MUX41X1 U1625 ( .IN1(reg13[3]), .IN3(reg15[3]), .IN2(reg14[3]), .IN4(
        reg16[3]), .S0(n1509), .S1(n1549), .Q(n1071) );
  MUX41X1 U1626 ( .IN1(reg9[3]), .IN3(reg11[3]), .IN2(reg10[3]), .IN4(reg12[3]), .S0(n1509), .S1(n1549), .Q(n1072) );
  MUX41X1 U1627 ( .IN1(reg5[3]), .IN3(reg7[3]), .IN2(reg6[3]), .IN4(reg8[3]), 
        .S0(n1509), .S1(n1549), .Q(n1073) );
  MUX41X1 U1628 ( .IN1(n1074), .IN3(n1072), .IN2(n1073), .IN4(n1071), .S0(
        n1488), .S1(n1494), .Q(n1075) );
  MUX21X1 U1629 ( .IN1(n1075), .IN2(n35), .S(n1484), .Q(rd_dataA[3]) );
  MUX41X1 U1630 ( .IN1(reg29[4]), .IN3(reg31[4]), .IN2(reg30[4]), .IN4(
        reg32[4]), .S0(n1509), .S1(n1549), .Q(n1076) );
  MUX41X1 U1631 ( .IN1(reg25[4]), .IN3(reg27[4]), .IN2(reg26[4]), .IN4(
        reg28[4]), .S0(n1509), .S1(n1549), .Q(n1077) );
  MUX41X1 U1632 ( .IN1(reg21[4]), .IN3(reg23[4]), .IN2(reg22[4]), .IN4(
        reg24[4]), .S0(n1509), .S1(n1549), .Q(n1078) );
  MUX41X1 U1633 ( .IN1(reg17[4]), .IN3(reg19[4]), .IN2(reg18[4]), .IN4(
        reg20[4]), .S0(n1509), .S1(n1549), .Q(n1079) );
  MUX41X1 U1634 ( .IN1(n1079), .IN3(n1077), .IN2(n1078), .IN4(n1076), .S0(
        n1488), .S1(n1494), .Q(n1080) );
  MUX41X1 U1635 ( .IN1(reg13[4]), .IN3(reg15[4]), .IN2(reg14[4]), .IN4(
        reg16[4]), .S0(n1509), .S1(n1549), .Q(n1081) );
  MUX41X1 U1636 ( .IN1(reg9[4]), .IN3(reg11[4]), .IN2(reg10[4]), .IN4(reg12[4]), .S0(n1509), .S1(n1549), .Q(n1082) );
  MUX41X1 U1637 ( .IN1(reg5[4]), .IN3(reg7[4]), .IN2(reg6[4]), .IN4(reg8[4]), 
        .S0(n1510), .S1(n1549), .Q(n1083) );
  MUX41X1 U1638 ( .IN1(n1084), .IN3(n1082), .IN2(n1083), .IN4(n1081), .S0(
        n1488), .S1(n1494), .Q(n1085) );
  MUX21X1 U1639 ( .IN1(n1085), .IN2(n1080), .S(n1484), .Q(rd_dataA[4]) );
  MUX41X1 U1640 ( .IN1(reg29[5]), .IN3(reg31[5]), .IN2(reg30[5]), .IN4(
        reg32[5]), .S0(n1510), .S1(n1549), .Q(n1086) );
  MUX41X1 U1641 ( .IN1(reg25[5]), .IN3(reg27[5]), .IN2(reg26[5]), .IN4(
        reg28[5]), .S0(n1510), .S1(n1549), .Q(n1087) );
  MUX41X1 U1642 ( .IN1(reg21[5]), .IN3(reg23[5]), .IN2(reg22[5]), .IN4(
        reg24[5]), .S0(n1510), .S1(n1550), .Q(n1088) );
  MUX41X1 U1643 ( .IN1(reg17[5]), .IN3(reg19[5]), .IN2(reg18[5]), .IN4(
        reg20[5]), .S0(n1510), .S1(n1550), .Q(n1089) );
  MUX41X1 U1644 ( .IN1(n1089), .IN3(n1087), .IN2(n1088), .IN4(n1086), .S0(
        n1488), .S1(n1494), .Q(n1090) );
  MUX41X1 U1645 ( .IN1(reg13[5]), .IN3(reg15[5]), .IN2(reg14[5]), .IN4(
        reg16[5]), .S0(n1510), .S1(n1550), .Q(n1091) );
  MUX41X1 U1646 ( .IN1(reg9[5]), .IN3(reg11[5]), .IN2(reg10[5]), .IN4(reg12[5]), .S0(n1510), .S1(n1550), .Q(n1092) );
  MUX41X1 U1647 ( .IN1(reg5[5]), .IN3(reg7[5]), .IN2(reg6[5]), .IN4(reg8[5]), 
        .S0(n1510), .S1(n1550), .Q(n1093) );
  MUX41X1 U1648 ( .IN1(n1094), .IN3(n1092), .IN2(n1093), .IN4(n1091), .S0(
        n1488), .S1(n1494), .Q(n1095) );
  MUX21X1 U1649 ( .IN1(n1095), .IN2(n1090), .S(n1484), .Q(rd_dataA[5]) );
  MUX41X1 U1650 ( .IN1(reg29[6]), .IN3(reg31[6]), .IN2(reg30[6]), .IN4(
        reg32[6]), .S0(n1510), .S1(n1550), .Q(n1096) );
  MUX41X1 U1651 ( .IN1(reg25[6]), .IN3(reg27[6]), .IN2(reg26[6]), .IN4(
        reg28[6]), .S0(n1510), .S1(n1550), .Q(n1097) );
  MUX41X1 U1652 ( .IN1(reg21[6]), .IN3(reg23[6]), .IN2(reg22[6]), .IN4(
        reg24[6]), .S0(n1510), .S1(n1550), .Q(n1098) );
  MUX41X1 U1653 ( .IN1(reg17[6]), .IN3(reg19[6]), .IN2(reg18[6]), .IN4(
        reg20[6]), .S0(n1510), .S1(n1550), .Q(n1099) );
  MUX41X1 U1654 ( .IN1(n1099), .IN3(n1097), .IN2(n1098), .IN4(n1096), .S0(
        n1488), .S1(n1494), .Q(n1100) );
  MUX41X1 U1655 ( .IN1(reg13[6]), .IN3(reg15[6]), .IN2(reg14[6]), .IN4(
        reg16[6]), .S0(n1510), .S1(n1550), .Q(n1101) );
  MUX41X1 U1656 ( .IN1(reg9[6]), .IN3(reg11[6]), .IN2(reg10[6]), .IN4(reg12[6]), .S0(n1510), .S1(n1550), .Q(n1102) );
  MUX41X1 U1657 ( .IN1(reg5[6]), .IN3(reg7[6]), .IN2(reg6[6]), .IN4(reg8[6]), 
        .S0(n1510), .S1(n1550), .Q(n1103) );
  MUX41X1 U1658 ( .IN1(n1104), .IN3(n1102), .IN2(n1103), .IN4(n1101), .S0(
        n1488), .S1(n1494), .Q(n1105) );
  MUX21X1 U1659 ( .IN1(n1105), .IN2(n1100), .S(n1484), .Q(rd_dataA[6]) );
  MUX41X1 U1660 ( .IN1(reg29[7]), .IN3(reg31[7]), .IN2(reg30[7]), .IN4(
        reg32[7]), .S0(n1511), .S1(n1551), .Q(n1106) );
  MUX41X1 U1661 ( .IN1(reg25[7]), .IN3(reg27[7]), .IN2(reg26[7]), .IN4(
        reg28[7]), .S0(n1511), .S1(n1551), .Q(n1107) );
  MUX41X1 U1662 ( .IN1(reg21[7]), .IN3(reg23[7]), .IN2(reg22[7]), .IN4(
        reg24[7]), .S0(n1511), .S1(n1551), .Q(n1108) );
  MUX41X1 U1663 ( .IN1(reg17[7]), .IN3(reg19[7]), .IN2(reg18[7]), .IN4(
        reg20[7]), .S0(n1511), .S1(n1551), .Q(n1109) );
  MUX41X1 U1664 ( .IN1(n1109), .IN3(n1107), .IN2(n1108), .IN4(n1106), .S0(
        n1488), .S1(n1494), .Q(n1110) );
  MUX41X1 U1665 ( .IN1(reg13[7]), .IN3(reg15[7]), .IN2(reg14[7]), .IN4(
        reg16[7]), .S0(n1511), .S1(n1551), .Q(n1111) );
  MUX41X1 U1666 ( .IN1(reg9[7]), .IN3(reg11[7]), .IN2(reg10[7]), .IN4(reg12[7]), .S0(n1511), .S1(n1551), .Q(n1112) );
  MUX41X1 U1667 ( .IN1(reg5[7]), .IN3(reg7[7]), .IN2(reg6[7]), .IN4(reg8[7]), 
        .S0(n1511), .S1(n1551), .Q(n1113) );
  MUX41X1 U1668 ( .IN1(n1114), .IN3(n1112), .IN2(n1113), .IN4(n1111), .S0(
        n1488), .S1(n1494), .Q(n1115) );
  MUX21X1 U1669 ( .IN1(n1115), .IN2(n1110), .S(n1484), .Q(rd_dataA[7]) );
  MUX41X1 U1670 ( .IN1(reg29[8]), .IN3(reg31[8]), .IN2(reg30[8]), .IN4(
        reg32[8]), .S0(n1511), .S1(n1551), .Q(n1116) );
  MUX41X1 U1671 ( .IN1(reg25[8]), .IN3(reg27[8]), .IN2(reg26[8]), .IN4(
        reg28[8]), .S0(n1511), .S1(n1551), .Q(n1117) );
  MUX41X1 U1672 ( .IN1(reg21[8]), .IN3(reg23[8]), .IN2(reg22[8]), .IN4(
        reg24[8]), .S0(n1511), .S1(n1551), .Q(n1118) );
  MUX41X1 U1673 ( .IN1(reg17[8]), .IN3(reg19[8]), .IN2(reg18[8]), .IN4(
        reg20[8]), .S0(n1511), .S1(n1551), .Q(n1119) );
  MUX41X1 U1674 ( .IN1(n1119), .IN3(n1117), .IN2(n1118), .IN4(n1116), .S0(
        n1489), .S1(n1495), .Q(n1120) );
  MUX41X1 U1675 ( .IN1(reg13[8]), .IN3(reg15[8]), .IN2(reg14[8]), .IN4(
        reg16[8]), .S0(n1511), .S1(n1551), .Q(n1121) );
  MUX41X1 U1676 ( .IN1(reg9[8]), .IN3(reg11[8]), .IN2(reg10[8]), .IN4(reg12[8]), .S0(n1511), .S1(n1552), .Q(n1122) );
  MUX41X1 U1677 ( .IN1(reg5[8]), .IN3(reg7[8]), .IN2(reg6[8]), .IN4(reg8[8]), 
        .S0(n1511), .S1(n1552), .Q(n1123) );
  MUX41X1 U1678 ( .IN1(n1124), .IN3(n1122), .IN2(n1123), .IN4(n1121), .S0(
        n1489), .S1(n1495), .Q(n1125) );
  MUX21X1 U1679 ( .IN1(n1125), .IN2(n1120), .S(n1485), .Q(rd_dataA[8]) );
  MUX41X1 U1680 ( .IN1(reg29[9]), .IN3(reg31[9]), .IN2(reg30[9]), .IN4(
        reg32[9]), .S0(n1511), .S1(n1552), .Q(n1126) );
  MUX41X1 U1681 ( .IN1(reg25[9]), .IN3(reg27[9]), .IN2(reg26[9]), .IN4(
        reg28[9]), .S0(n1512), .S1(n1552), .Q(n1127) );
  MUX41X1 U1682 ( .IN1(reg21[9]), .IN3(reg23[9]), .IN2(reg22[9]), .IN4(
        reg24[9]), .S0(n1512), .S1(n1552), .Q(n1128) );
  MUX41X1 U1683 ( .IN1(reg17[9]), .IN3(reg19[9]), .IN2(reg18[9]), .IN4(
        reg20[9]), .S0(n1512), .S1(n1552), .Q(n1129) );
  MUX41X1 U1684 ( .IN1(n1129), .IN3(n1127), .IN2(n1128), .IN4(n1126), .S0(
        n1489), .S1(n1495), .Q(n1130) );
  MUX41X1 U1685 ( .IN1(reg13[9]), .IN3(reg15[9]), .IN2(reg14[9]), .IN4(
        reg16[9]), .S0(n1512), .S1(n1552), .Q(n1131) );
  MUX41X1 U1686 ( .IN1(reg9[9]), .IN3(reg11[9]), .IN2(reg10[9]), .IN4(reg12[9]), .S0(n1512), .S1(n1552), .Q(n1132) );
  MUX41X1 U1687 ( .IN1(reg5[9]), .IN3(reg7[9]), .IN2(reg6[9]), .IN4(reg8[9]), 
        .S0(n1512), .S1(n1552), .Q(n1133) );
  MUX41X1 U1688 ( .IN1(n1134), .IN3(n1132), .IN2(n1133), .IN4(n1131), .S0(
        n1489), .S1(n1495), .Q(n1135) );
  MUX21X1 U1689 ( .IN1(n1135), .IN2(n1130), .S(n1485), .Q(rd_dataA[9]) );
  MUX41X1 U1690 ( .IN1(reg29[10]), .IN3(reg31[10]), .IN2(reg30[10]), .IN4(
        reg32[10]), .S0(n1512), .S1(n1552), .Q(n1136) );
  MUX41X1 U1691 ( .IN1(reg25[10]), .IN3(reg27[10]), .IN2(reg26[10]), .IN4(
        reg28[10]), .S0(n1512), .S1(n1552), .Q(n1137) );
  MUX41X1 U1692 ( .IN1(reg21[10]), .IN3(reg23[10]), .IN2(reg22[10]), .IN4(
        reg24[10]), .S0(n1512), .S1(n1552), .Q(n1138) );
  MUX41X1 U1693 ( .IN1(reg17[10]), .IN3(reg19[10]), .IN2(reg18[10]), .IN4(
        reg20[10]), .S0(n1512), .S1(n1553), .Q(n1139) );
  MUX41X1 U1694 ( .IN1(n1139), .IN3(n1137), .IN2(n1138), .IN4(n1136), .S0(
        n1489), .S1(n1495), .Q(n1140) );
  MUX41X1 U1695 ( .IN1(reg13[10]), .IN3(reg15[10]), .IN2(reg14[10]), .IN4(
        reg16[10]), .S0(n1512), .S1(n1553), .Q(n1141) );
  MUX41X1 U1696 ( .IN1(reg9[10]), .IN3(reg11[10]), .IN2(reg10[10]), .IN4(
        reg12[10]), .S0(n1512), .S1(n1553), .Q(n1142) );
  MUX41X1 U1697 ( .IN1(reg5[10]), .IN3(reg7[10]), .IN2(reg6[10]), .IN4(
        reg8[10]), .S0(n1512), .S1(n1553), .Q(n1143) );
  MUX41X1 U1698 ( .IN1(n1144), .IN3(n1142), .IN2(n1143), .IN4(n1141), .S0(
        n1489), .S1(n1495), .Q(n1145) );
  MUX21X1 U1699 ( .IN1(n1145), .IN2(n1140), .S(n1485), .Q(rd_dataA[10]) );
  MUX41X1 U1700 ( .IN1(reg29[11]), .IN3(reg31[11]), .IN2(reg30[11]), .IN4(
        reg32[11]), .S0(n1512), .S1(n1553), .Q(n1146) );
  MUX41X1 U1701 ( .IN1(reg25[11]), .IN3(reg27[11]), .IN2(reg26[11]), .IN4(
        reg28[11]), .S0(n1513), .S1(n1553), .Q(n1147) );
  MUX41X1 U1702 ( .IN1(reg21[11]), .IN3(reg23[11]), .IN2(reg22[11]), .IN4(
        reg24[11]), .S0(n1513), .S1(n1553), .Q(n1148) );
  MUX41X1 U1703 ( .IN1(reg17[11]), .IN3(reg19[11]), .IN2(reg18[11]), .IN4(
        reg20[11]), .S0(n1513), .S1(n1553), .Q(n1149) );
  MUX41X1 U1704 ( .IN1(n1149), .IN3(n1147), .IN2(n1148), .IN4(n1146), .S0(
        n1489), .S1(n1495), .Q(n1150) );
  MUX41X1 U1705 ( .IN1(reg13[11]), .IN3(reg15[11]), .IN2(reg14[11]), .IN4(
        reg16[11]), .S0(n1513), .S1(n1553), .Q(n1151) );
  MUX41X1 U1706 ( .IN1(reg9[11]), .IN3(reg11[11]), .IN2(reg10[11]), .IN4(
        reg12[11]), .S0(n1513), .S1(n1553), .Q(n1152) );
  MUX41X1 U1707 ( .IN1(reg5[11]), .IN3(reg7[11]), .IN2(reg6[11]), .IN4(
        reg8[11]), .S0(n1513), .S1(n1553), .Q(n1153) );
  MUX41X1 U1708 ( .IN1(n1154), .IN3(n1152), .IN2(n1153), .IN4(n1151), .S0(
        n1489), .S1(n1495), .Q(n1155) );
  MUX21X1 U1709 ( .IN1(n1155), .IN2(n1150), .S(n1485), .Q(rd_dataA[11]) );
  MUX41X1 U1710 ( .IN1(reg29[12]), .IN3(reg31[12]), .IN2(reg30[12]), .IN4(
        reg32[12]), .S0(n1513), .S1(n1554), .Q(n1156) );
  MUX41X1 U1711 ( .IN1(reg25[12]), .IN3(reg27[12]), .IN2(reg26[12]), .IN4(
        reg28[12]), .S0(n1513), .S1(n1554), .Q(n1157) );
  MUX41X1 U1712 ( .IN1(reg21[12]), .IN3(reg23[12]), .IN2(reg22[12]), .IN4(
        reg24[12]), .S0(n1513), .S1(n1554), .Q(n1158) );
  MUX41X1 U1713 ( .IN1(reg17[12]), .IN3(reg19[12]), .IN2(reg18[12]), .IN4(
        reg20[12]), .S0(n1513), .S1(n1554), .Q(n1159) );
  MUX41X1 U1714 ( .IN1(n1159), .IN3(n1157), .IN2(n1158), .IN4(n1156), .S0(
        n1489), .S1(n1495), .Q(n1160) );
  MUX41X1 U1715 ( .IN1(reg13[12]), .IN3(reg15[12]), .IN2(reg14[12]), .IN4(
        reg16[12]), .S0(n1513), .S1(n1554), .Q(n1161) );
  MUX41X1 U1716 ( .IN1(reg9[12]), .IN3(reg11[12]), .IN2(reg10[12]), .IN4(
        reg12[12]), .S0(n1513), .S1(n1554), .Q(n1162) );
  MUX41X1 U1717 ( .IN1(reg5[12]), .IN3(reg7[12]), .IN2(reg6[12]), .IN4(
        reg8[12]), .S0(n1513), .S1(n1554), .Q(n1163) );
  MUX41X1 U1718 ( .IN1(n1164), .IN3(n1162), .IN2(n1163), .IN4(n1161), .S0(
        n1489), .S1(n1495), .Q(n1165) );
  MUX21X1 U1719 ( .IN1(n1165), .IN2(n1160), .S(n1485), .Q(rd_dataA[12]) );
  MUX41X1 U1720 ( .IN1(reg29[13]), .IN3(reg31[13]), .IN2(reg30[13]), .IN4(
        reg32[13]), .S0(n1513), .S1(n1554), .Q(n1166) );
  MUX41X1 U1721 ( .IN1(reg25[13]), .IN3(reg27[13]), .IN2(reg26[13]), .IN4(
        reg28[13]), .S0(n1513), .S1(n1554), .Q(n1167) );
  MUX41X1 U1722 ( .IN1(reg21[13]), .IN3(reg23[13]), .IN2(reg22[13]), .IN4(
        reg24[13]), .S0(n1514), .S1(n1554), .Q(n1168) );
  MUX41X1 U1723 ( .IN1(reg17[13]), .IN3(reg19[13]), .IN2(reg18[13]), .IN4(
        reg20[13]), .S0(n1514), .S1(n1554), .Q(n1169) );
  MUX41X1 U1724 ( .IN1(n1169), .IN3(n1167), .IN2(n1168), .IN4(n1166), .S0(
        n1489), .S1(n1495), .Q(n1170) );
  MUX41X1 U1725 ( .IN1(reg13[13]), .IN3(reg15[13]), .IN2(reg14[13]), .IN4(
        reg16[13]), .S0(n1514), .S1(n1554), .Q(n1171) );
  MUX41X1 U1726 ( .IN1(reg9[13]), .IN3(reg11[13]), .IN2(reg10[13]), .IN4(
        reg12[13]), .S0(n1514), .S1(n1555), .Q(n1172) );
  MUX41X1 U1727 ( .IN1(reg5[13]), .IN3(reg7[13]), .IN2(reg6[13]), .IN4(
        reg8[13]), .S0(n1514), .S1(n1556), .Q(n1173) );
  MUX41X1 U1728 ( .IN1(n1174), .IN3(n1172), .IN2(n1173), .IN4(n1171), .S0(
        n1489), .S1(n1495), .Q(n1175) );
  MUX21X1 U1729 ( .IN1(n1175), .IN2(n1170), .S(n1485), .Q(rd_dataA[13]) );
  MUX41X1 U1730 ( .IN1(reg29[14]), .IN3(reg31[14]), .IN2(reg30[14]), .IN4(
        reg32[14]), .S0(n1514), .S1(n1542), .Q(n1176) );
  MUX41X1 U1731 ( .IN1(reg25[14]), .IN3(reg27[14]), .IN2(reg26[14]), .IN4(
        reg28[14]), .S0(n1514), .S1(n1543), .Q(n1177) );
  MUX41X1 U1732 ( .IN1(reg21[14]), .IN3(reg23[14]), .IN2(reg22[14]), .IN4(
        reg24[14]), .S0(n1514), .S1(n1545), .Q(n1178) );
  MUX41X1 U1733 ( .IN1(reg17[14]), .IN3(reg19[14]), .IN2(reg18[14]), .IN4(
        reg20[14]), .S0(n1514), .S1(n1541), .Q(n1179) );
  MUX41X1 U1734 ( .IN1(n1179), .IN3(n1177), .IN2(n1178), .IN4(n1176), .S0(
        n1490), .S1(n1496), .Q(n1180) );
  MUX41X1 U1735 ( .IN1(reg13[14]), .IN3(reg15[14]), .IN2(reg14[14]), .IN4(
        reg16[14]), .S0(n1514), .S1(n1546), .Q(n1181) );
  MUX41X1 U1736 ( .IN1(reg9[14]), .IN3(reg11[14]), .IN2(reg10[14]), .IN4(
        reg12[14]), .S0(n1514), .S1(n1544), .Q(n1182) );
  MUX41X1 U1737 ( .IN1(reg5[14]), .IN3(reg7[14]), .IN2(reg6[14]), .IN4(
        reg8[14]), .S0(n1514), .S1(n1538), .Q(n1183) );
  MUX41X1 U1738 ( .IN1(n1184), .IN3(n1182), .IN2(n1183), .IN4(n1181), .S0(
        n1490), .S1(n1496), .Q(n1185) );
  MUX21X1 U1739 ( .IN1(n1185), .IN2(n1180), .S(n1485), .Q(rd_dataA[14]) );
  MUX41X1 U1740 ( .IN1(reg29[15]), .IN3(reg31[15]), .IN2(reg30[15]), .IN4(
        reg32[15]), .S0(n1515), .S1(n1545), .Q(n1186) );
  MUX41X1 U1741 ( .IN1(reg25[15]), .IN3(reg27[15]), .IN2(reg26[15]), .IN4(
        reg28[15]), .S0(n1515), .S1(n1546), .Q(n1187) );
  MUX41X1 U1742 ( .IN1(reg21[15]), .IN3(reg23[15]), .IN2(reg22[15]), .IN4(
        reg24[15]), .S0(n1514), .S1(n1544), .Q(n1188) );
  MUX41X1 U1743 ( .IN1(reg17[15]), .IN3(reg19[15]), .IN2(reg18[15]), .IN4(
        reg20[15]), .S0(n1515), .S1(n1555), .Q(n1189) );
  MUX41X1 U1744 ( .IN1(n1189), .IN3(n1187), .IN2(n1188), .IN4(n1186), .S0(
        n1490), .S1(n1496), .Q(n1190) );
  MUX41X1 U1745 ( .IN1(reg13[15]), .IN3(reg15[15]), .IN2(reg14[15]), .IN4(
        reg16[15]), .S0(n1515), .S1(n1555), .Q(n1191) );
  MUX41X1 U1746 ( .IN1(reg9[15]), .IN3(reg11[15]), .IN2(reg10[15]), .IN4(
        reg12[15]), .S0(n1514), .S1(n1555), .Q(n1192) );
  MUX41X1 U1747 ( .IN1(reg5[15]), .IN3(reg7[15]), .IN2(reg6[15]), .IN4(
        reg8[15]), .S0(n1515), .S1(n1555), .Q(n1193) );
  MUX41X1 U1748 ( .IN1(n1194), .IN3(n1192), .IN2(n1193), .IN4(n1191), .S0(
        n1490), .S1(n1496), .Q(n1195) );
  MUX21X1 U1749 ( .IN1(n1195), .IN2(n1190), .S(n1485), .Q(rd_dataA[15]) );
  MUX41X1 U1750 ( .IN1(reg29[16]), .IN3(reg31[16]), .IN2(reg30[16]), .IN4(
        reg32[16]), .S0(n1515), .S1(n1555), .Q(n1196) );
  MUX41X1 U1751 ( .IN1(reg25[16]), .IN3(reg27[16]), .IN2(reg26[16]), .IN4(
        reg28[16]), .S0(n1515), .S1(n1555), .Q(n1197) );
  MUX41X1 U1752 ( .IN1(reg21[16]), .IN3(reg23[16]), .IN2(reg22[16]), .IN4(
        reg24[16]), .S0(n1515), .S1(n1555), .Q(n1198) );
  MUX41X1 U1753 ( .IN1(reg17[16]), .IN3(reg19[16]), .IN2(reg18[16]), .IN4(
        reg20[16]), .S0(n1515), .S1(n1555), .Q(n1199) );
  MUX41X1 U1754 ( .IN1(n1199), .IN3(n1197), .IN2(n1198), .IN4(n1196), .S0(
        n1490), .S1(n1496), .Q(n1200) );
  MUX41X1 U1755 ( .IN1(reg13[16]), .IN3(reg15[16]), .IN2(reg14[16]), .IN4(
        reg16[16]), .S0(n1515), .S1(n1555), .Q(n1201) );
  MUX41X1 U1756 ( .IN1(reg9[16]), .IN3(reg11[16]), .IN2(reg10[16]), .IN4(
        reg12[16]), .S0(n1515), .S1(n1555), .Q(n1202) );
  MUX41X1 U1757 ( .IN1(reg5[16]), .IN3(reg7[16]), .IN2(reg6[16]), .IN4(
        reg8[16]), .S0(n1514), .S1(n1555), .Q(n1203) );
  MUX41X1 U1758 ( .IN1(n1204), .IN3(n1202), .IN2(n1203), .IN4(n1201), .S0(
        n1490), .S1(n1496), .Q(n1205) );
  MUX21X1 U1759 ( .IN1(n1205), .IN2(n1200), .S(n1485), .Q(rd_dataA[16]) );
  MUX41X1 U1760 ( .IN1(reg29[17]), .IN3(reg31[17]), .IN2(reg30[17]), .IN4(
        reg32[17]), .S0(n1515), .S1(n1555), .Q(n1206) );
  MUX41X1 U1761 ( .IN1(reg25[17]), .IN3(reg27[17]), .IN2(reg26[17]), .IN4(
        reg28[17]), .S0(n1515), .S1(n1556), .Q(n1207) );
  MUX41X1 U1762 ( .IN1(reg21[17]), .IN3(reg23[17]), .IN2(reg22[17]), .IN4(
        reg24[17]), .S0(n1516), .S1(n1556), .Q(n1208) );
  MUX41X1 U1763 ( .IN1(reg17[17]), .IN3(reg19[17]), .IN2(reg18[17]), .IN4(
        reg20[17]), .S0(n1515), .S1(n1556), .Q(n1209) );
  MUX41X1 U1764 ( .IN1(n1209), .IN3(n1207), .IN2(n1208), .IN4(n1206), .S0(
        n1490), .S1(n1496), .Q(n1210) );
  MUX41X1 U1765 ( .IN1(reg13[17]), .IN3(reg15[17]), .IN2(reg14[17]), .IN4(
        reg16[17]), .S0(n1516), .S1(n1556), .Q(n1211) );
  MUX41X1 U1766 ( .IN1(reg9[17]), .IN3(reg11[17]), .IN2(reg10[17]), .IN4(
        reg12[17]), .S0(n1516), .S1(n1556), .Q(n1212) );
  MUX41X1 U1767 ( .IN1(reg5[17]), .IN3(reg7[17]), .IN2(reg6[17]), .IN4(
        reg8[17]), .S0(n1515), .S1(n1556), .Q(n1213) );
  MUX41X1 U1768 ( .IN1(n1214), .IN3(n1212), .IN2(n1213), .IN4(n1211), .S0(
        n1490), .S1(n1496), .Q(n1215) );
  MUX21X1 U1769 ( .IN1(n1215), .IN2(n1210), .S(n1485), .Q(rd_dataA[17]) );
  MUX41X1 U1770 ( .IN1(reg29[18]), .IN3(reg31[18]), .IN2(reg30[18]), .IN4(
        reg32[18]), .S0(n1516), .S1(n1556), .Q(n1216) );
  MUX41X1 U1771 ( .IN1(reg25[18]), .IN3(reg27[18]), .IN2(reg26[18]), .IN4(
        reg28[18]), .S0(n1512), .S1(n1556), .Q(n1217) );
  MUX41X1 U1772 ( .IN1(reg21[18]), .IN3(reg23[18]), .IN2(reg22[18]), .IN4(
        reg24[18]), .S0(n1501), .S1(n1556), .Q(n1218) );
  MUX41X1 U1773 ( .IN1(reg17[18]), .IN3(reg19[18]), .IN2(reg18[18]), .IN4(
        reg20[18]), .S0(n1501), .S1(n1556), .Q(n1219) );
  MUX41X1 U1774 ( .IN1(n1219), .IN3(n1217), .IN2(n1218), .IN4(n1216), .S0(
        n1490), .S1(n1496), .Q(n1220) );
  MUX41X1 U1775 ( .IN1(reg13[18]), .IN3(reg15[18]), .IN2(reg14[18]), .IN4(
        reg16[18]), .S0(n1501), .S1(n1556), .Q(n1221) );
  MUX41X1 U1776 ( .IN1(reg9[18]), .IN3(reg11[18]), .IN2(reg10[18]), .IN4(
        reg12[18]), .S0(n1501), .S1(n1556), .Q(n1222) );
  MUX41X1 U1777 ( .IN1(reg5[18]), .IN3(reg7[18]), .IN2(reg6[18]), .IN4(
        reg8[18]), .S0(n1501), .S1(n1557), .Q(n1223) );
  MUX41X1 U1778 ( .IN1(n1224), .IN3(n1222), .IN2(n1223), .IN4(n1221), .S0(
        n1490), .S1(n1496), .Q(n1225) );
  MUX21X1 U1779 ( .IN1(n1225), .IN2(n1220), .S(n1485), .Q(rd_dataA[18]) );
  MUX41X1 U1780 ( .IN1(reg29[19]), .IN3(reg31[19]), .IN2(reg30[19]), .IN4(
        reg32[19]), .S0(n1501), .S1(n1557), .Q(n1226) );
  MUX41X1 U1781 ( .IN1(reg25[19]), .IN3(reg27[19]), .IN2(reg26[19]), .IN4(
        reg28[19]), .S0(n1501), .S1(n1557), .Q(n1227) );
  MUX41X1 U1782 ( .IN1(reg21[19]), .IN3(reg23[19]), .IN2(reg22[19]), .IN4(
        reg24[19]), .S0(n1501), .S1(n1557), .Q(n1228) );
  MUX41X1 U1783 ( .IN1(reg17[19]), .IN3(reg19[19]), .IN2(reg18[19]), .IN4(
        reg20[19]), .S0(n1501), .S1(n1557), .Q(n1229) );
  MUX41X1 U1784 ( .IN1(n1229), .IN3(n1227), .IN2(n1228), .IN4(n1226), .S0(
        n1490), .S1(n1496), .Q(n1230) );
  MUX41X1 U1785 ( .IN1(reg13[19]), .IN3(reg15[19]), .IN2(reg14[19]), .IN4(
        reg16[19]), .S0(n1502), .S1(n1557), .Q(n1231) );
  MUX41X1 U1786 ( .IN1(reg9[19]), .IN3(reg11[19]), .IN2(reg10[19]), .IN4(
        reg12[19]), .S0(n1502), .S1(n1557), .Q(n1232) );
  MUX41X1 U1787 ( .IN1(reg5[19]), .IN3(reg7[19]), .IN2(reg6[19]), .IN4(
        reg8[19]), .S0(n1502), .S1(n1557), .Q(n1233) );
  MUX41X1 U1788 ( .IN1(n1234), .IN3(n1232), .IN2(n1233), .IN4(n1231), .S0(
        n1490), .S1(n1496), .Q(n1235) );
  MUX21X1 U1789 ( .IN1(n1235), .IN2(n1230), .S(n1485), .Q(rd_dataA[19]) );
  MUX41X1 U1790 ( .IN1(reg29[20]), .IN3(reg31[20]), .IN2(reg30[20]), .IN4(
        reg32[20]), .S0(n1502), .S1(n1557), .Q(n1236) );
  MUX41X1 U1791 ( .IN1(reg25[20]), .IN3(reg27[20]), .IN2(reg26[20]), .IN4(
        reg28[20]), .S0(n1502), .S1(n1557), .Q(n1237) );
  MUX41X1 U1792 ( .IN1(reg21[20]), .IN3(reg23[20]), .IN2(reg22[20]), .IN4(
        reg24[20]), .S0(n1502), .S1(n1557), .Q(n1238) );
  MUX41X1 U1793 ( .IN1(reg17[20]), .IN3(reg19[20]), .IN2(reg18[20]), .IN4(
        reg20[20]), .S0(n1502), .S1(n1553), .Q(n1239) );
  MUX41X1 U1794 ( .IN1(n1239), .IN3(n1237), .IN2(n1238), .IN4(n1236), .S0(
        n1491), .S1(n1497), .Q(n1240) );
  MUX41X1 U1795 ( .IN1(reg13[20]), .IN3(reg15[20]), .IN2(reg14[20]), .IN4(
        reg16[20]), .S0(n1504), .S1(n1543), .Q(n1241) );
  MUX41X1 U1796 ( .IN1(reg9[20]), .IN3(reg11[20]), .IN2(reg10[20]), .IN4(
        reg12[20]), .S0(n1502), .S1(n1540), .Q(n1242) );
  MUX41X1 U1797 ( .IN1(reg5[20]), .IN3(reg7[20]), .IN2(reg6[20]), .IN4(
        reg8[20]), .S0(n1502), .S1(n1540), .Q(n1243) );
  MUX41X1 U1798 ( .IN1(n1244), .IN3(n1242), .IN2(n1243), .IN4(n1241), .S0(
        n1491), .S1(n1497), .Q(n1245) );
  MUX21X1 U1799 ( .IN1(n1245), .IN2(n1240), .S(n1486), .Q(rd_dataA[20]) );
  MUX41X1 U1800 ( .IN1(reg29[21]), .IN3(reg31[21]), .IN2(reg30[21]), .IN4(
        reg32[21]), .S0(n1502), .S1(n1540), .Q(n1246) );
  MUX41X1 U1801 ( .IN1(reg25[21]), .IN3(reg27[21]), .IN2(reg26[21]), .IN4(
        reg28[21]), .S0(n1502), .S1(n1540), .Q(n1247) );
  MUX41X1 U1802 ( .IN1(reg21[21]), .IN3(reg23[21]), .IN2(reg22[21]), .IN4(
        reg24[21]), .S0(n1502), .S1(n1540), .Q(n1248) );
  MUX41X1 U1803 ( .IN1(reg17[21]), .IN3(reg19[21]), .IN2(reg18[21]), .IN4(
        reg20[21]), .S0(n1502), .S1(n1540), .Q(n1249) );
  MUX41X1 U1804 ( .IN1(n1249), .IN3(n1247), .IN2(n1248), .IN4(n1246), .S0(
        n1491), .S1(n1497), .Q(n1250) );
  MUX41X1 U1805 ( .IN1(reg13[21]), .IN3(reg15[21]), .IN2(reg14[21]), .IN4(
        reg16[21]), .S0(n1502), .S1(n1540), .Q(n1251) );
  MUX41X1 U1806 ( .IN1(reg9[21]), .IN3(reg11[21]), .IN2(reg10[21]), .IN4(
        reg12[21]), .S0(n1503), .S1(n1541), .Q(n1252) );
  MUX41X1 U1807 ( .IN1(reg5[21]), .IN3(reg7[21]), .IN2(reg6[21]), .IN4(
        reg8[21]), .S0(n1503), .S1(n1541), .Q(n1253) );
  MUX41X1 U1808 ( .IN1(n1254), .IN3(n1252), .IN2(n1253), .IN4(n1251), .S0(
        n1491), .S1(n1497), .Q(n1255) );
  MUX21X1 U1809 ( .IN1(n1255), .IN2(n1250), .S(n1486), .Q(rd_dataA[21]) );
  MUX41X1 U1810 ( .IN1(reg29[22]), .IN3(reg31[22]), .IN2(reg30[22]), .IN4(
        reg32[22]), .S0(n1503), .S1(n1541), .Q(n1256) );
  MUX41X1 U1811 ( .IN1(reg25[22]), .IN3(reg27[22]), .IN2(reg26[22]), .IN4(
        reg28[22]), .S0(n1503), .S1(n1541), .Q(n1257) );
  MUX41X1 U1812 ( .IN1(reg21[22]), .IN3(reg23[22]), .IN2(reg22[22]), .IN4(
        reg24[22]), .S0(n1503), .S1(n1541), .Q(n1258) );
  MUX41X1 U1813 ( .IN1(reg17[22]), .IN3(reg19[22]), .IN2(reg18[22]), .IN4(
        reg20[22]), .S0(n1503), .S1(n1541), .Q(n1259) );
  MUX41X1 U1814 ( .IN1(n1259), .IN3(n1257), .IN2(n1258), .IN4(n1256), .S0(
        n1491), .S1(n1497), .Q(n1260) );
  MUX41X1 U1815 ( .IN1(reg13[22]), .IN3(reg15[22]), .IN2(reg14[22]), .IN4(
        reg16[22]), .S0(n1503), .S1(n1541), .Q(n1261) );
  MUX41X1 U1816 ( .IN1(reg9[22]), .IN3(reg11[22]), .IN2(reg10[22]), .IN4(
        reg12[22]), .S0(n1503), .S1(n1541), .Q(n1262) );
  MUX41X1 U1817 ( .IN1(reg5[22]), .IN3(reg7[22]), .IN2(reg6[22]), .IN4(
        reg8[22]), .S0(n1503), .S1(n1541), .Q(n1263) );
  MUX41X1 U1818 ( .IN1(n1264), .IN3(n1262), .IN2(n1263), .IN4(n1261), .S0(
        n1491), .S1(n1497), .Q(n1265) );
  MUX21X1 U1819 ( .IN1(n1265), .IN2(n1260), .S(n1486), .Q(rd_dataA[22]) );
  MUX41X1 U1820 ( .IN1(reg29[23]), .IN3(reg31[23]), .IN2(reg30[23]), .IN4(
        reg32[23]), .S0(n1503), .S1(n1541), .Q(n1266) );
  MUX41X1 U1821 ( .IN1(reg25[23]), .IN3(reg27[23]), .IN2(reg26[23]), .IN4(
        reg28[23]), .S0(n1503), .S1(n1541), .Q(n1267) );
  MUX41X1 U1822 ( .IN1(reg21[23]), .IN3(reg23[23]), .IN2(reg22[23]), .IN4(
        reg24[23]), .S0(n1503), .S1(n1541), .Q(n1268) );
  MUX41X1 U1823 ( .IN1(reg17[23]), .IN3(reg19[23]), .IN2(reg18[23]), .IN4(
        reg20[23]), .S0(n1503), .S1(n1542), .Q(n1269) );
  MUX41X1 U1824 ( .IN1(n1269), .IN3(n1267), .IN2(n1268), .IN4(n1266), .S0(
        n1491), .S1(n1497), .Q(n1270) );
  MUX41X1 U1825 ( .IN1(reg13[23]), .IN3(reg15[23]), .IN2(reg14[23]), .IN4(
        reg16[23]), .S0(n1503), .S1(n1542), .Q(n1271) );
  MUX41X1 U1826 ( .IN1(reg9[23]), .IN3(reg11[23]), .IN2(reg10[23]), .IN4(
        reg12[23]), .S0(n1503), .S1(n1542), .Q(n1272) );
  MUX41X1 U1827 ( .IN1(reg5[23]), .IN3(reg7[23]), .IN2(reg6[23]), .IN4(
        reg8[23]), .S0(n1504), .S1(n1542), .Q(n1273) );
  MUX41X1 U1828 ( .IN1(n1274), .IN3(n1272), .IN2(n1273), .IN4(n1271), .S0(
        n1491), .S1(n1497), .Q(n1275) );
  MUX21X1 U1829 ( .IN1(n1275), .IN2(n1270), .S(n1486), .Q(rd_dataA[23]) );
  MUX41X1 U1830 ( .IN1(reg29[24]), .IN3(reg31[24]), .IN2(reg30[24]), .IN4(
        reg32[24]), .S0(n1504), .S1(n1542), .Q(n1276) );
  MUX41X1 U1831 ( .IN1(reg25[24]), .IN3(reg27[24]), .IN2(reg26[24]), .IN4(
        reg28[24]), .S0(n1504), .S1(n1542), .Q(n1277) );
  MUX41X1 U1832 ( .IN1(reg21[24]), .IN3(reg23[24]), .IN2(reg22[24]), .IN4(
        reg24[24]), .S0(n1504), .S1(n1542), .Q(n1278) );
  MUX41X1 U1833 ( .IN1(reg17[24]), .IN3(reg19[24]), .IN2(reg18[24]), .IN4(
        reg20[24]), .S0(n1504), .S1(n1542), .Q(n1279) );
  MUX41X1 U1834 ( .IN1(n1279), .IN3(n1277), .IN2(n1278), .IN4(n1276), .S0(
        n1491), .S1(n1497), .Q(n1280) );
  MUX41X1 U1835 ( .IN1(reg13[24]), .IN3(reg15[24]), .IN2(reg14[24]), .IN4(
        reg16[24]), .S0(n1504), .S1(n1542), .Q(n1281) );
  MUX41X1 U1836 ( .IN1(reg9[24]), .IN3(reg11[24]), .IN2(reg10[24]), .IN4(
        reg12[24]), .S0(n1504), .S1(n1542), .Q(n1282) );
  MUX41X1 U1837 ( .IN1(reg5[24]), .IN3(reg7[24]), .IN2(reg6[24]), .IN4(
        reg8[24]), .S0(n1504), .S1(n1542), .Q(n1283) );
  MUX41X1 U1838 ( .IN1(n1284), .IN3(n1282), .IN2(n1283), .IN4(n1281), .S0(
        n1491), .S1(n1497), .Q(n1285) );
  MUX21X1 U1839 ( .IN1(n1285), .IN2(n1280), .S(n1486), .Q(rd_dataA[24]) );
  MUX41X1 U1840 ( .IN1(reg29[25]), .IN3(reg31[25]), .IN2(reg30[25]), .IN4(
        reg32[25]), .S0(n1504), .S1(n1542), .Q(n1286) );
  MUX41X1 U1841 ( .IN1(reg25[25]), .IN3(reg27[25]), .IN2(reg26[25]), .IN4(
        reg28[25]), .S0(n1504), .S1(n1543), .Q(n1287) );
  MUX41X1 U1842 ( .IN1(reg21[25]), .IN3(reg23[25]), .IN2(reg22[25]), .IN4(
        reg24[25]), .S0(n1504), .S1(n1543), .Q(n1288) );
  MUX41X1 U1843 ( .IN1(reg17[25]), .IN3(reg19[25]), .IN2(reg18[25]), .IN4(
        reg20[25]), .S0(n1504), .S1(n1543), .Q(n1289) );
  MUX41X1 U1844 ( .IN1(n1289), .IN3(n1287), .IN2(n1288), .IN4(n1286), .S0(
        n1491), .S1(n1497), .Q(n1290) );
  MUX41X1 U1845 ( .IN1(reg13[25]), .IN3(reg15[25]), .IN2(reg14[25]), .IN4(
        reg16[25]), .S0(n1504), .S1(n1543), .Q(n1291) );
  MUX41X1 U1846 ( .IN1(reg9[25]), .IN3(reg11[25]), .IN2(reg10[25]), .IN4(
        reg12[25]), .S0(n1504), .S1(n1543), .Q(n1292) );
  MUX41X1 U1847 ( .IN1(reg5[25]), .IN3(reg7[25]), .IN2(reg6[25]), .IN4(
        reg8[25]), .S0(n1505), .S1(n1543), .Q(n1293) );
  MUX41X1 U1848 ( .IN1(n1294), .IN3(n1292), .IN2(n1293), .IN4(n1291), .S0(
        n1491), .S1(n1497), .Q(n1295) );
  MUX21X1 U1849 ( .IN1(n1295), .IN2(n1290), .S(n1486), .Q(rd_dataA[25]) );
  MUX41X1 U1850 ( .IN1(reg29[26]), .IN3(reg31[26]), .IN2(reg30[26]), .IN4(
        reg32[26]), .S0(n1505), .S1(n1543), .Q(n1296) );
  MUX41X1 U1851 ( .IN1(reg25[26]), .IN3(reg27[26]), .IN2(reg26[26]), .IN4(
        reg28[26]), .S0(n1505), .S1(n1543), .Q(n1297) );
  MUX41X1 U1852 ( .IN1(reg21[26]), .IN3(reg23[26]), .IN2(reg22[26]), .IN4(
        reg24[26]), .S0(n1505), .S1(n1543), .Q(n1298) );
  MUX41X1 U1853 ( .IN1(reg17[26]), .IN3(reg19[26]), .IN2(reg18[26]), .IN4(
        reg20[26]), .S0(n1505), .S1(n1543), .Q(n1299) );
  MUX41X1 U1854 ( .IN1(n1299), .IN3(n1297), .IN2(n1298), .IN4(n1296), .S0(
        n1492), .S1(n1498), .Q(n1300) );
  MUX41X1 U1855 ( .IN1(reg13[26]), .IN3(reg15[26]), .IN2(reg14[26]), .IN4(
        reg16[26]), .S0(n1505), .S1(n1543), .Q(n1301) );
  MUX41X1 U1856 ( .IN1(reg9[26]), .IN3(reg11[26]), .IN2(reg10[26]), .IN4(
        reg12[26]), .S0(n1505), .S1(n1544), .Q(n1302) );
  MUX41X1 U1857 ( .IN1(reg5[26]), .IN3(reg7[26]), .IN2(reg6[26]), .IN4(
        reg8[26]), .S0(n1505), .S1(n1544), .Q(n1303) );
  MUX41X1 U1858 ( .IN1(n1304), .IN3(n1302), .IN2(n1303), .IN4(n1301), .S0(
        n1492), .S1(n1498), .Q(n1305) );
  MUX21X1 U1859 ( .IN1(n1305), .IN2(n1300), .S(n1486), .Q(rd_dataA[26]) );
  MUX41X1 U1860 ( .IN1(reg29[27]), .IN3(reg31[27]), .IN2(reg30[27]), .IN4(
        reg32[27]), .S0(n1505), .S1(n1544), .Q(n1306) );
  MUX41X1 U1861 ( .IN1(reg25[27]), .IN3(reg27[27]), .IN2(reg26[27]), .IN4(
        reg28[27]), .S0(n1505), .S1(n1544), .Q(n1307) );
  MUX41X1 U1862 ( .IN1(reg21[27]), .IN3(reg23[27]), .IN2(reg22[27]), .IN4(
        reg24[27]), .S0(n1505), .S1(n1544), .Q(n1308) );
  MUX41X1 U1863 ( .IN1(reg17[27]), .IN3(reg19[27]), .IN2(reg18[27]), .IN4(
        reg20[27]), .S0(n1505), .S1(n1544), .Q(n1309) );
  MUX41X1 U1864 ( .IN1(n1309), .IN3(n1307), .IN2(n1308), .IN4(n1306), .S0(
        n1492), .S1(n1498), .Q(n1310) );
  MUX41X1 U1865 ( .IN1(reg13[27]), .IN3(reg15[27]), .IN2(reg14[27]), .IN4(
        reg16[27]), .S0(n1505), .S1(n1544), .Q(n1311) );
  MUX41X1 U1866 ( .IN1(reg9[27]), .IN3(reg11[27]), .IN2(reg10[27]), .IN4(
        reg12[27]), .S0(n1505), .S1(n1544), .Q(n1312) );
  MUX41X1 U1867 ( .IN1(reg5[27]), .IN3(reg7[27]), .IN2(reg6[27]), .IN4(
        reg8[27]), .S0(n1505), .S1(n1544), .Q(n1313) );
  MUX41X1 U1868 ( .IN1(n1314), .IN3(n1312), .IN2(n1313), .IN4(n1311), .S0(
        n1492), .S1(n1498), .Q(n1315) );
  MUX21X1 U1869 ( .IN1(n1315), .IN2(n1310), .S(n1486), .Q(rd_dataA[27]) );
  MUX41X1 U1870 ( .IN1(reg29[28]), .IN3(reg31[28]), .IN2(reg30[28]), .IN4(
        reg32[28]), .S0(n1506), .S1(n1544), .Q(n1316) );
  MUX41X1 U1871 ( .IN1(reg25[28]), .IN3(reg27[28]), .IN2(reg26[28]), .IN4(
        reg28[28]), .S0(n1506), .S1(n1544), .Q(n1317) );
  MUX41X1 U1872 ( .IN1(reg21[28]), .IN3(reg23[28]), .IN2(reg22[28]), .IN4(
        reg24[28]), .S0(n1506), .S1(n1544), .Q(n1318) );
  MUX41X1 U1873 ( .IN1(reg17[28]), .IN3(reg19[28]), .IN2(reg18[28]), .IN4(
        reg20[28]), .S0(n1506), .S1(n1545), .Q(n1319) );
  MUX41X1 U1874 ( .IN1(n1319), .IN3(n1317), .IN2(n1318), .IN4(n1316), .S0(
        n1492), .S1(n1498), .Q(n1320) );
  MUX41X1 U1875 ( .IN1(reg13[28]), .IN3(reg15[28]), .IN2(reg14[28]), .IN4(
        reg16[28]), .S0(n1506), .S1(n1545), .Q(n1321) );
  MUX41X1 U1876 ( .IN1(reg9[28]), .IN3(reg11[28]), .IN2(reg10[28]), .IN4(
        reg12[28]), .S0(n1506), .S1(n1545), .Q(n1322) );
  MUX41X1 U1877 ( .IN1(reg5[28]), .IN3(reg7[28]), .IN2(reg6[28]), .IN4(
        reg8[28]), .S0(n1506), .S1(n1545), .Q(n1323) );
  MUX41X1 U1878 ( .IN1(n1324), .IN3(n1322), .IN2(n1323), .IN4(n1321), .S0(
        n1492), .S1(n1498), .Q(n1325) );
  MUX21X1 U1879 ( .IN1(n1325), .IN2(n1320), .S(n1486), .Q(rd_dataA[28]) );
  MUX41X1 U1880 ( .IN1(reg29[29]), .IN3(reg31[29]), .IN2(reg30[29]), .IN4(
        reg32[29]), .S0(n1506), .S1(n1545), .Q(n1326) );
  MUX41X1 U1881 ( .IN1(reg25[29]), .IN3(reg27[29]), .IN2(reg26[29]), .IN4(
        reg28[29]), .S0(n1506), .S1(n1545), .Q(n1327) );
  MUX41X1 U1882 ( .IN1(reg21[29]), .IN3(reg23[29]), .IN2(reg22[29]), .IN4(
        reg24[29]), .S0(n1506), .S1(n1545), .Q(n1328) );
  MUX41X1 U1883 ( .IN1(reg17[29]), .IN3(reg19[29]), .IN2(reg18[29]), .IN4(
        reg20[29]), .S0(n1506), .S1(n1545), .Q(n1329) );
  MUX41X1 U1884 ( .IN1(n1329), .IN3(n1327), .IN2(n1328), .IN4(n1326), .S0(
        n1492), .S1(n1498), .Q(n1330) );
  MUX41X1 U1885 ( .IN1(reg13[29]), .IN3(reg15[29]), .IN2(reg14[29]), .IN4(
        reg16[29]), .S0(n1506), .S1(n1545), .Q(n1331) );
  MUX41X1 U1886 ( .IN1(reg9[29]), .IN3(reg11[29]), .IN2(reg10[29]), .IN4(
        reg12[29]), .S0(n1506), .S1(n1545), .Q(n1332) );
  MUX41X1 U1887 ( .IN1(reg5[29]), .IN3(reg7[29]), .IN2(reg6[29]), .IN4(
        reg8[29]), .S0(n1506), .S1(n1545), .Q(n1333) );
  MUX41X1 U1888 ( .IN1(n1334), .IN3(n1332), .IN2(n1333), .IN4(n1331), .S0(
        n1492), .S1(n1498), .Q(n1335) );
  MUX21X1 U1889 ( .IN1(n1335), .IN2(n1330), .S(n1486), .Q(rd_dataA[29]) );
  MUX41X1 U1890 ( .IN1(reg29[30]), .IN3(reg31[30]), .IN2(reg30[30]), .IN4(
        reg32[30]), .S0(n1506), .S1(n1545), .Q(n1336) );
  MUX41X1 U1891 ( .IN1(reg25[30]), .IN3(reg27[30]), .IN2(reg26[30]), .IN4(
        reg28[30]), .S0(n1507), .S1(n1546), .Q(n1337) );
  MUX41X1 U1892 ( .IN1(reg21[30]), .IN3(reg23[30]), .IN2(reg22[30]), .IN4(
        reg24[30]), .S0(n1507), .S1(n1546), .Q(n1338) );
  MUX41X1 U1893 ( .IN1(reg17[30]), .IN3(reg19[30]), .IN2(reg18[30]), .IN4(
        reg20[30]), .S0(n1507), .S1(n1546), .Q(n1339) );
  MUX41X1 U1894 ( .IN1(n1339), .IN3(n1337), .IN2(n1338), .IN4(n1336), .S0(
        n1492), .S1(n1498), .Q(n1340) );
  MUX41X1 U1895 ( .IN1(reg13[30]), .IN3(reg15[30]), .IN2(reg14[30]), .IN4(
        reg16[30]), .S0(n1507), .S1(n1546), .Q(n1341) );
  MUX41X1 U1896 ( .IN1(reg9[30]), .IN3(reg11[30]), .IN2(reg10[30]), .IN4(
        reg12[30]), .S0(n1507), .S1(n1546), .Q(n1342) );
  MUX41X1 U1897 ( .IN1(reg5[30]), .IN3(reg7[30]), .IN2(reg6[30]), .IN4(
        reg8[30]), .S0(n1507), .S1(n1546), .Q(n1343) );
  MUX41X1 U1898 ( .IN1(n1344), .IN3(n1342), .IN2(n1343), .IN4(n1341), .S0(
        n1492), .S1(n1498), .Q(n1345) );
  MUX21X1 U1899 ( .IN1(n1345), .IN2(n1340), .S(n1486), .Q(rd_dataA[30]) );
  MUX41X1 U1900 ( .IN1(reg29[31]), .IN3(reg31[31]), .IN2(reg30[31]), .IN4(
        reg32[31]), .S0(n1507), .S1(n1546), .Q(n1346) );
  MUX41X1 U1901 ( .IN1(reg25[31]), .IN3(reg27[31]), .IN2(reg26[31]), .IN4(
        reg28[31]), .S0(n1507), .S1(n1546), .Q(n1347) );
  MUX41X1 U1902 ( .IN1(reg21[31]), .IN3(reg23[31]), .IN2(reg22[31]), .IN4(
        reg24[31]), .S0(n1507), .S1(n1546), .Q(n1348) );
  MUX41X1 U1903 ( .IN1(reg17[31]), .IN3(reg19[31]), .IN2(reg18[31]), .IN4(
        reg20[31]), .S0(n1507), .S1(n1546), .Q(n1349) );
  MUX41X1 U1904 ( .IN1(n1349), .IN3(n1347), .IN2(n1348), .IN4(n1346), .S0(
        n1492), .S1(n1498), .Q(n1350) );
  MUX41X1 U1905 ( .IN1(reg13[31]), .IN3(reg15[31]), .IN2(reg14[31]), .IN4(
        reg16[31]), .S0(n1507), .S1(n1546), .Q(n1351) );
  MUX41X1 U1906 ( .IN1(reg9[31]), .IN3(reg11[31]), .IN2(reg10[31]), .IN4(
        reg12[31]), .S0(n1507), .S1(n1546), .Q(n1352) );
  MUX41X1 U1907 ( .IN1(reg5[31]), .IN3(reg7[31]), .IN2(reg6[31]), .IN4(
        reg8[31]), .S0(n1507), .S1(n1547), .Q(n1353) );
  MUX41X1 U1908 ( .IN1(n1354), .IN3(n1352), .IN2(n1353), .IN4(n1351), .S0(
        n1492), .S1(n1498), .Q(n1355) );
  MUX21X1 U1909 ( .IN1(n1355), .IN2(n1350), .S(n1486), .Q(rd_dataA[31]) );
  MUX21X1 U1910 ( .IN1(n1356), .IN2(n1357), .S(n1516), .Q(n1359) );
  NAND3X0 U1911 ( .IN1(reg4[31]), .IN2(n1501), .IN3(n1536), .QN(n1358) );
  MUX21X1 U1912 ( .IN1(n1360), .IN2(n1361), .S(n1517), .Q(n1363) );
  NAND3X0 U1913 ( .IN1(reg4[30]), .IN2(n1501), .IN3(n1536), .QN(n1362) );
  MUX21X1 U1914 ( .IN1(n1364), .IN2(n1365), .S(n1516), .Q(n1367) );
  NAND3X0 U1915 ( .IN1(reg4[29]), .IN2(n1501), .IN3(n1536), .QN(n1366) );
  MUX21X1 U1916 ( .IN1(n1368), .IN2(n1369), .S(n1516), .Q(n1371) );
  NAND3X0 U1917 ( .IN1(reg4[28]), .IN2(n1501), .IN3(n1537), .QN(n1370) );
  MUX21X1 U1918 ( .IN1(n1372), .IN2(n1373), .S(n1517), .Q(n1375) );
  NAND3X0 U1919 ( .IN1(reg4[27]), .IN2(n1501), .IN3(n1537), .QN(n1374) );
  MUX21X1 U1920 ( .IN1(n1376), .IN2(n1377), .S(n1516), .Q(n1379) );
  NAND3X0 U1921 ( .IN1(reg4[26]), .IN2(n1501), .IN3(n1537), .QN(n1378) );
  MUX21X1 U1922 ( .IN1(n1380), .IN2(n1381), .S(n1516), .Q(n1383) );
  NAND3X0 U1923 ( .IN1(reg4[25]), .IN2(n1501), .IN3(n1537), .QN(n1382) );
  MUX21X1 U1924 ( .IN1(n1384), .IN2(n1385), .S(n1517), .Q(n1387) );
  NAND3X0 U1925 ( .IN1(reg4[24]), .IN2(n1500), .IN3(n1537), .QN(n1386) );
  MUX21X1 U1926 ( .IN1(n1388), .IN2(n1389), .S(n1516), .Q(n1391) );
  NAND3X0 U1927 ( .IN1(reg4[23]), .IN2(n1500), .IN3(n1537), .QN(n1390) );
  MUX21X1 U1928 ( .IN1(n1392), .IN2(n1393), .S(n1516), .Q(n1395) );
  NAND3X0 U1929 ( .IN1(reg4[22]), .IN2(n1500), .IN3(n1537), .QN(n1394) );
  MUX21X1 U1930 ( .IN1(n1396), .IN2(n1397), .S(n1517), .Q(n1399) );
  NAND3X0 U1931 ( .IN1(reg4[21]), .IN2(n1500), .IN3(n1537), .QN(n1398) );
  MUX21X1 U1932 ( .IN1(n1400), .IN2(n1401), .S(n1516), .Q(n1403) );
  NAND3X0 U1933 ( .IN1(reg4[20]), .IN2(n1500), .IN3(n1537), .QN(n1402) );
  MUX21X1 U1934 ( .IN1(n1404), .IN2(n1405), .S(n1517), .Q(n1407) );
  NAND3X0 U1935 ( .IN1(reg4[19]), .IN2(n1500), .IN3(n1537), .QN(n1406) );
  MUX21X1 U1936 ( .IN1(n1408), .IN2(n1409), .S(n1517), .Q(n1411) );
  NAND3X0 U1937 ( .IN1(reg4[18]), .IN2(n1500), .IN3(n1537), .QN(n1410) );
  MUX21X1 U1938 ( .IN1(n1412), .IN2(n1413), .S(n1517), .Q(n1415) );
  NAND3X0 U1939 ( .IN1(reg4[17]), .IN2(n1500), .IN3(n1537), .QN(n1414) );
  MUX21X1 U1940 ( .IN1(n1416), .IN2(n1417), .S(n1517), .Q(n1419) );
  NAND3X0 U1941 ( .IN1(reg4[16]), .IN2(n1500), .IN3(n1537), .QN(n1418) );
  MUX21X1 U1942 ( .IN1(n1420), .IN2(n1421), .S(n1518), .Q(n1423) );
  NAND3X0 U1943 ( .IN1(reg4[15]), .IN2(n1500), .IN3(n1537), .QN(n1422) );
  MUX21X1 U1944 ( .IN1(n1424), .IN2(n1425), .S(n1517), .Q(n1427) );
  NAND3X0 U1945 ( .IN1(reg4[14]), .IN2(n1500), .IN3(n1537), .QN(n1426) );
  MUX21X1 U1946 ( .IN1(n1428), .IN2(n1429), .S(n1517), .Q(n1431) );
  NAND3X0 U1947 ( .IN1(reg4[13]), .IN2(n1500), .IN3(n1537), .QN(n1430) );
  MUX21X1 U1948 ( .IN1(n1432), .IN2(n1433), .S(n1518), .Q(n1435) );
  NAND3X0 U1949 ( .IN1(reg4[12]), .IN2(n1500), .IN3(n1537), .QN(n1434) );
  MUX21X1 U1950 ( .IN1(n1436), .IN2(n1437), .S(n1517), .Q(n1439) );
  NAND3X0 U1951 ( .IN1(reg4[11]), .IN2(n1500), .IN3(n1537), .QN(n1438) );
  MUX21X1 U1952 ( .IN1(n1440), .IN2(n1441), .S(n1517), .Q(n1443) );
  NAND3X0 U1953 ( .IN1(reg4[10]), .IN2(n1500), .IN3(n1537), .QN(n1442) );
  MUX21X1 U1954 ( .IN1(n1444), .IN2(n1445), .S(n1518), .Q(n1447) );
  NAND3X0 U1955 ( .IN1(reg4[9]), .IN2(n1500), .IN3(n1537), .QN(n1446) );
  MUX21X1 U1956 ( .IN1(n1448), .IN2(n1449), .S(n1518), .Q(n1451) );
  NAND3X0 U1957 ( .IN1(reg4[8]), .IN2(n1500), .IN3(n1537), .QN(n1450) );
  MUX21X1 U1958 ( .IN1(n1452), .IN2(n1453), .S(n1518), .Q(n1455) );
  NAND3X0 U1959 ( .IN1(reg4[7]), .IN2(n1500), .IN3(n1537), .QN(n1454) );
  MUX21X1 U1960 ( .IN1(n1456), .IN2(n1457), .S(n1518), .Q(n1459) );
  NAND3X0 U1961 ( .IN1(reg4[6]), .IN2(n1499), .IN3(n1536), .QN(n1458) );
  MUX21X1 U1962 ( .IN1(n1460), .IN2(n1461), .S(n1518), .Q(n1463) );
  NAND3X0 U1963 ( .IN1(reg4[5]), .IN2(n1499), .IN3(n1537), .QN(n1462) );
  MUX21X1 U1964 ( .IN1(n1464), .IN2(n1465), .S(n1518), .Q(n1467) );
  NAND3X0 U1965 ( .IN1(reg4[4]), .IN2(n1499), .IN3(n1536), .QN(n1466) );
  MUX21X1 U1966 ( .IN1(n1468), .IN2(n1469), .S(n1518), .Q(n1471) );
  NAND3X0 U1967 ( .IN1(reg4[3]), .IN2(n1499), .IN3(n1536), .QN(n1470) );
  MUX21X1 U1968 ( .IN1(n1472), .IN2(n1473), .S(n1518), .Q(n1475) );
  NAND3X0 U1969 ( .IN1(reg4[2]), .IN2(n1499), .IN3(n1536), .QN(n1474) );
  MUX21X1 U1970 ( .IN1(n1476), .IN2(n1477), .S(n1518), .Q(n1479) );
  NAND3X0 U1971 ( .IN1(reg4[1]), .IN2(n1499), .IN3(n1536), .QN(n1478) );
  MUX21X1 U1972 ( .IN1(n1480), .IN2(n1481), .S(n1518), .Q(n1483) );
  NAND3X0 U1973 ( .IN1(reg4[0]), .IN2(n1499), .IN3(n1537), .QN(n1482) );
  INVX0 U1974 ( .INP(N11), .ZN(n1521) );
  INVX0 U1975 ( .INP(n1522), .ZN(n1536) );
  INVX0 U1976 ( .INP(n1523), .ZN(n1538) );
  INVX0 U1977 ( .INP(n1523), .ZN(n1539) );
  INVX0 U1978 ( .INP(n1523), .ZN(n1540) );
  INVX0 U1979 ( .INP(n1523), .ZN(n1541) );
  INVX0 U1980 ( .INP(n1523), .ZN(n1542) );
  INVX0 U1981 ( .INP(n1523), .ZN(n1543) );
  INVX0 U1982 ( .INP(n1523), .ZN(n1544) );
  INVX0 U1983 ( .INP(n1523), .ZN(n1545) );
  INVX0 U1984 ( .INP(n1523), .ZN(n1546) );
  INVX0 U1985 ( .INP(n1524), .ZN(n1547) );
  INVX0 U1986 ( .INP(n1524), .ZN(n1548) );
  INVX0 U1987 ( .INP(n1524), .ZN(n1549) );
  INVX0 U1988 ( .INP(n1524), .ZN(n1550) );
  INVX0 U1989 ( .INP(n1524), .ZN(n1551) );
  INVX0 U1990 ( .INP(n1524), .ZN(n1552) );
  INVX0 U1991 ( .INP(n1524), .ZN(n1553) );
  INVX0 U1992 ( .INP(n1524), .ZN(n1554) );
  MUX41X1 U1993 ( .IN1(reg29[0]), .IN3(reg31[0]), .IN2(reg30[0]), .IN4(
        reg32[0]), .S0(n2024), .S1(n2062), .Q(n1558) );
  MUX41X1 U1994 ( .IN1(reg25[0]), .IN3(reg27[0]), .IN2(reg26[0]), .IN4(
        reg28[0]), .S0(n2038), .S1(n2079), .Q(n1559) );
  MUX41X1 U1995 ( .IN1(reg21[0]), .IN3(reg23[0]), .IN2(reg22[0]), .IN4(
        reg24[0]), .S0(n2029), .S1(n2069), .Q(n1560) );
  MUX41X1 U1996 ( .IN1(reg17[0]), .IN3(reg19[0]), .IN2(reg18[0]), .IN4(
        reg20[0]), .S0(n2029), .S1(n2069), .Q(n1561) );
  MUX41X1 U1997 ( .IN1(n1561), .IN3(n1559), .IN2(n1560), .IN4(n1558), .S0(
        n2009), .S1(n2015), .Q(n1562) );
  MUX41X1 U1998 ( .IN1(reg13[0]), .IN3(reg15[0]), .IN2(reg14[0]), .IN4(
        reg16[0]), .S0(n2030), .S1(n2069), .Q(n1563) );
  MUX41X1 U1999 ( .IN1(reg9[0]), .IN3(reg11[0]), .IN2(reg10[0]), .IN4(reg12[0]), .S0(n2030), .S1(n2069), .Q(n1564) );
  MUX41X1 U2000 ( .IN1(reg5[0]), .IN3(reg7[0]), .IN2(reg6[0]), .IN4(reg8[0]), 
        .S0(n2030), .S1(n2069), .Q(n1565) );
  MUX41X1 U2001 ( .IN1(n1566), .IN3(n1564), .IN2(n1565), .IN4(n1563), .S0(
        n2009), .S1(n2015), .Q(n1567) );
  MUX21X1 U2002 ( .IN1(n1567), .IN2(n1562), .S(n2006), .Q(rd_dataB[0]) );
  MUX41X1 U2003 ( .IN1(reg29[1]), .IN3(reg31[1]), .IN2(reg30[1]), .IN4(
        reg32[1]), .S0(n2030), .S1(n2069), .Q(n1568) );
  MUX41X1 U2004 ( .IN1(reg25[1]), .IN3(reg27[1]), .IN2(reg26[1]), .IN4(
        reg28[1]), .S0(n2030), .S1(n2069), .Q(n1569) );
  MUX41X1 U2005 ( .IN1(reg21[1]), .IN3(reg23[1]), .IN2(reg22[1]), .IN4(
        reg24[1]), .S0(n2030), .S1(n2069), .Q(n1570) );
  MUX41X1 U2006 ( .IN1(reg17[1]), .IN3(reg19[1]), .IN2(reg18[1]), .IN4(
        reg20[1]), .S0(n2030), .S1(n2069), .Q(n1571) );
  MUX41X1 U2007 ( .IN1(n1571), .IN3(n1569), .IN2(n1570), .IN4(n1568), .S0(
        n2009), .S1(n2015), .Q(n1572) );
  MUX41X1 U2008 ( .IN1(reg13[1]), .IN3(reg15[1]), .IN2(reg14[1]), .IN4(
        reg16[1]), .S0(n2030), .S1(n2069), .Q(n1573) );
  MUX41X1 U2009 ( .IN1(reg9[1]), .IN3(reg11[1]), .IN2(reg10[1]), .IN4(reg12[1]), .S0(n2030), .S1(n2069), .Q(n1574) );
  MUX41X1 U2010 ( .IN1(reg5[1]), .IN3(reg7[1]), .IN2(reg6[1]), .IN4(reg8[1]), 
        .S0(n2030), .S1(n2070), .Q(n1575) );
  MUX41X1 U2011 ( .IN1(n1576), .IN3(n1574), .IN2(n1575), .IN4(n1573), .S0(
        n2009), .S1(n2015), .Q(n1577) );
  MUX21X1 U2012 ( .IN1(n1577), .IN2(n1572), .S(n2006), .Q(rd_dataB[1]) );
  MUX41X1 U2013 ( .IN1(reg29[2]), .IN3(reg31[2]), .IN2(reg30[2]), .IN4(
        reg32[2]), .S0(n2030), .S1(n2070), .Q(n1578) );
  MUX41X1 U2014 ( .IN1(reg25[2]), .IN3(reg27[2]), .IN2(reg26[2]), .IN4(
        reg28[2]), .S0(n2030), .S1(n2070), .Q(n1579) );
  MUX41X1 U2015 ( .IN1(reg21[2]), .IN3(reg23[2]), .IN2(reg22[2]), .IN4(
        reg24[2]), .S0(n2030), .S1(n2070), .Q(n1580) );
  MUX41X1 U2016 ( .IN1(reg17[2]), .IN3(reg19[2]), .IN2(reg18[2]), .IN4(
        reg20[2]), .S0(n2030), .S1(n2070), .Q(n1581) );
  MUX41X1 U2017 ( .IN1(n1581), .IN3(n1579), .IN2(n1580), .IN4(n1578), .S0(
        n2010), .S1(n2016), .Q(n1582) );
  MUX41X1 U2018 ( .IN1(reg13[2]), .IN3(reg15[2]), .IN2(reg14[2]), .IN4(
        reg16[2]), .S0(n2030), .S1(n2070), .Q(n1583) );
  MUX41X1 U2019 ( .IN1(reg9[2]), .IN3(reg11[2]), .IN2(reg10[2]), .IN4(reg12[2]), .S0(n2031), .S1(n2070), .Q(n1584) );
  MUX41X1 U2020 ( .IN1(reg5[2]), .IN3(reg7[2]), .IN2(reg6[2]), .IN4(reg8[2]), 
        .S0(n2031), .S1(n2070), .Q(n1585) );
  MUX41X1 U2021 ( .IN1(n1586), .IN3(n1584), .IN2(n1585), .IN4(n1583), .S0(
        n2010), .S1(n2016), .Q(n1587) );
  MUX21X1 U2022 ( .IN1(n1587), .IN2(n1582), .S(n2006), .Q(rd_dataB[2]) );
  MUX41X1 U2023 ( .IN1(reg29[3]), .IN3(reg31[3]), .IN2(reg30[3]), .IN4(
        reg32[3]), .S0(n2031), .S1(n2070), .Q(n1588) );
  MUX41X1 U2024 ( .IN1(reg25[3]), .IN3(reg27[3]), .IN2(reg26[3]), .IN4(
        reg28[3]), .S0(n2031), .S1(n2070), .Q(n1589) );
  MUX41X1 U2025 ( .IN1(reg21[3]), .IN3(reg23[3]), .IN2(reg22[3]), .IN4(
        reg24[3]), .S0(n2031), .S1(n2070), .Q(n1590) );
  MUX41X1 U2026 ( .IN1(reg17[3]), .IN3(reg19[3]), .IN2(reg18[3]), .IN4(
        reg20[3]), .S0(n2031), .S1(n2070), .Q(n1591) );
  MUX41X1 U2027 ( .IN1(n1591), .IN3(n1589), .IN2(n1590), .IN4(n1588), .S0(
        n2010), .S1(n2016), .Q(n1592) );
  MUX41X1 U2028 ( .IN1(reg13[3]), .IN3(reg15[3]), .IN2(reg14[3]), .IN4(
        reg16[3]), .S0(n2031), .S1(n2071), .Q(n1593) );
  MUX41X1 U2029 ( .IN1(reg9[3]), .IN3(reg11[3]), .IN2(reg10[3]), .IN4(reg12[3]), .S0(n2031), .S1(n2071), .Q(n1594) );
  MUX41X1 U2030 ( .IN1(reg5[3]), .IN3(reg7[3]), .IN2(reg6[3]), .IN4(reg8[3]), 
        .S0(n2031), .S1(n2071), .Q(n1595) );
  MUX41X1 U2031 ( .IN1(n1596), .IN3(n1594), .IN2(n1595), .IN4(n1593), .S0(
        n2010), .S1(n2016), .Q(n1597) );
  MUX21X1 U2032 ( .IN1(n1597), .IN2(n1592), .S(n2006), .Q(rd_dataB[3]) );
  MUX41X1 U2033 ( .IN1(reg29[4]), .IN3(reg31[4]), .IN2(reg30[4]), .IN4(
        reg32[4]), .S0(n2031), .S1(n2071), .Q(n1598) );
  MUX41X1 U2034 ( .IN1(reg25[4]), .IN3(reg27[4]), .IN2(reg26[4]), .IN4(
        reg28[4]), .S0(n2031), .S1(n2071), .Q(n1599) );
  MUX41X1 U2035 ( .IN1(reg21[4]), .IN3(reg23[4]), .IN2(reg22[4]), .IN4(
        reg24[4]), .S0(n2031), .S1(n2071), .Q(n1600) );
  MUX41X1 U2036 ( .IN1(reg17[4]), .IN3(reg19[4]), .IN2(reg18[4]), .IN4(
        reg20[4]), .S0(n2031), .S1(n2071), .Q(n1601) );
  MUX41X1 U2037 ( .IN1(n1601), .IN3(n1599), .IN2(n1600), .IN4(n1598), .S0(
        n2010), .S1(n2016), .Q(n1602) );
  MUX41X1 U2038 ( .IN1(reg13[4]), .IN3(reg15[4]), .IN2(reg14[4]), .IN4(
        reg16[4]), .S0(n2031), .S1(n2071), .Q(n1603) );
  MUX41X1 U2039 ( .IN1(reg9[4]), .IN3(reg11[4]), .IN2(reg10[4]), .IN4(reg12[4]), .S0(n2031), .S1(n2071), .Q(n1604) );
  MUX41X1 U2040 ( .IN1(reg5[4]), .IN3(reg7[4]), .IN2(reg6[4]), .IN4(reg8[4]), 
        .S0(n2032), .S1(n2071), .Q(n1605) );
  MUX41X1 U2041 ( .IN1(n1606), .IN3(n1604), .IN2(n1605), .IN4(n1603), .S0(
        n2010), .S1(n2016), .Q(n1607) );
  MUX21X1 U2042 ( .IN1(n1607), .IN2(n1602), .S(n2006), .Q(rd_dataB[4]) );
  MUX41X1 U2043 ( .IN1(reg29[5]), .IN3(reg31[5]), .IN2(reg30[5]), .IN4(
        reg32[5]), .S0(n2032), .S1(n2071), .Q(n1608) );
  MUX41X1 U2044 ( .IN1(reg25[5]), .IN3(reg27[5]), .IN2(reg26[5]), .IN4(
        reg28[5]), .S0(n2032), .S1(n2071), .Q(n1609) );
  MUX41X1 U2045 ( .IN1(reg21[5]), .IN3(reg23[5]), .IN2(reg22[5]), .IN4(
        reg24[5]), .S0(n2032), .S1(n2072), .Q(n1610) );
  MUX41X1 U2046 ( .IN1(reg17[5]), .IN3(reg19[5]), .IN2(reg18[5]), .IN4(
        reg20[5]), .S0(n2032), .S1(n2072), .Q(n1611) );
  MUX41X1 U2047 ( .IN1(n1611), .IN3(n1609), .IN2(n1610), .IN4(n1608), .S0(
        n2010), .S1(n2016), .Q(n1612) );
  MUX41X1 U2048 ( .IN1(reg13[5]), .IN3(reg15[5]), .IN2(reg14[5]), .IN4(
        reg16[5]), .S0(n2032), .S1(n2072), .Q(n1613) );
  MUX41X1 U2049 ( .IN1(reg9[5]), .IN3(reg11[5]), .IN2(reg10[5]), .IN4(reg12[5]), .S0(n2032), .S1(n2072), .Q(n1614) );
  MUX41X1 U2050 ( .IN1(reg5[5]), .IN3(reg7[5]), .IN2(reg6[5]), .IN4(reg8[5]), 
        .S0(n2032), .S1(n2072), .Q(n1615) );
  MUX41X1 U2051 ( .IN1(n1616), .IN3(n1614), .IN2(n1615), .IN4(n1613), .S0(
        n2010), .S1(n2016), .Q(n1617) );
  MUX21X1 U2052 ( .IN1(n1617), .IN2(n1612), .S(n2006), .Q(rd_dataB[5]) );
  MUX41X1 U2053 ( .IN1(reg29[6]), .IN3(reg31[6]), .IN2(reg30[6]), .IN4(
        reg32[6]), .S0(n2032), .S1(n2072), .Q(n1618) );
  MUX41X1 U2054 ( .IN1(reg25[6]), .IN3(reg27[6]), .IN2(reg26[6]), .IN4(
        reg28[6]), .S0(n2032), .S1(n2072), .Q(n1619) );
  MUX41X1 U2055 ( .IN1(reg21[6]), .IN3(reg23[6]), .IN2(reg22[6]), .IN4(
        reg24[6]), .S0(n2032), .S1(n2072), .Q(n1620) );
  MUX41X1 U2056 ( .IN1(reg17[6]), .IN3(reg19[6]), .IN2(reg18[6]), .IN4(
        reg20[6]), .S0(n2032), .S1(n2072), .Q(n1621) );
  MUX41X1 U2057 ( .IN1(n1621), .IN3(n1619), .IN2(n1620), .IN4(n1618), .S0(
        n2010), .S1(n2016), .Q(n1622) );
  MUX41X1 U2058 ( .IN1(reg13[6]), .IN3(reg15[6]), .IN2(reg14[6]), .IN4(
        reg16[6]), .S0(n2032), .S1(n2072), .Q(n1623) );
  MUX41X1 U2059 ( .IN1(reg9[6]), .IN3(reg11[6]), .IN2(reg10[6]), .IN4(reg12[6]), .S0(n2032), .S1(n2072), .Q(n1624) );
  MUX41X1 U2060 ( .IN1(reg5[6]), .IN3(reg7[6]), .IN2(reg6[6]), .IN4(reg8[6]), 
        .S0(n2032), .S1(n2072), .Q(n1625) );
  MUX41X1 U2061 ( .IN1(n1626), .IN3(n1624), .IN2(n1625), .IN4(n1623), .S0(
        n2010), .S1(n2016), .Q(n1627) );
  MUX21X1 U2062 ( .IN1(n1627), .IN2(n1622), .S(n2006), .Q(rd_dataB[6]) );
  MUX41X1 U2063 ( .IN1(reg29[7]), .IN3(reg31[7]), .IN2(reg30[7]), .IN4(
        reg32[7]), .S0(n2033), .S1(n2073), .Q(n1628) );
  MUX41X1 U2064 ( .IN1(reg25[7]), .IN3(reg27[7]), .IN2(reg26[7]), .IN4(
        reg28[7]), .S0(n2033), .S1(n2073), .Q(n1629) );
  MUX41X1 U2065 ( .IN1(reg21[7]), .IN3(reg23[7]), .IN2(reg22[7]), .IN4(
        reg24[7]), .S0(n2033), .S1(n2073), .Q(n1630) );
  MUX41X1 U2066 ( .IN1(reg17[7]), .IN3(reg19[7]), .IN2(reg18[7]), .IN4(
        reg20[7]), .S0(n2033), .S1(n2073), .Q(n1631) );
  MUX41X1 U2067 ( .IN1(n1631), .IN3(n1629), .IN2(n1630), .IN4(n1628), .S0(
        n2010), .S1(n2016), .Q(n1632) );
  MUX41X1 U2068 ( .IN1(reg13[7]), .IN3(reg15[7]), .IN2(reg14[7]), .IN4(
        reg16[7]), .S0(n2033), .S1(n2073), .Q(n1633) );
  MUX41X1 U2069 ( .IN1(reg9[7]), .IN3(reg11[7]), .IN2(reg10[7]), .IN4(reg12[7]), .S0(n2033), .S1(n2073), .Q(n1634) );
  MUX41X1 U2070 ( .IN1(reg5[7]), .IN3(reg7[7]), .IN2(reg6[7]), .IN4(reg8[7]), 
        .S0(n2033), .S1(n2073), .Q(n1635) );
  MUX41X1 U2071 ( .IN1(n1636), .IN3(n1634), .IN2(n1635), .IN4(n1633), .S0(
        n2010), .S1(n2016), .Q(n1637) );
  MUX21X1 U2072 ( .IN1(n1637), .IN2(n1632), .S(n2006), .Q(rd_dataB[7]) );
  MUX41X1 U2073 ( .IN1(reg29[8]), .IN3(reg31[8]), .IN2(reg30[8]), .IN4(
        reg32[8]), .S0(n2033), .S1(n2073), .Q(n1638) );
  MUX41X1 U2074 ( .IN1(reg25[8]), .IN3(reg27[8]), .IN2(reg26[8]), .IN4(
        reg28[8]), .S0(n2033), .S1(n2073), .Q(n1639) );
  MUX41X1 U2075 ( .IN1(reg21[8]), .IN3(reg23[8]), .IN2(reg22[8]), .IN4(
        reg24[8]), .S0(n2033), .S1(n2073), .Q(n1640) );
  MUX41X1 U2076 ( .IN1(reg17[8]), .IN3(reg19[8]), .IN2(reg18[8]), .IN4(
        reg20[8]), .S0(n2033), .S1(n2073), .Q(n1641) );
  MUX41X1 U2077 ( .IN1(n1641), .IN3(n1639), .IN2(n1640), .IN4(n1638), .S0(
        n2011), .S1(n2017), .Q(n1642) );
  MUX41X1 U2078 ( .IN1(reg13[8]), .IN3(reg15[8]), .IN2(reg14[8]), .IN4(
        reg16[8]), .S0(n2033), .S1(n2073), .Q(n1643) );
  MUX41X1 U2079 ( .IN1(reg9[8]), .IN3(reg11[8]), .IN2(reg10[8]), .IN4(reg12[8]), .S0(n2033), .S1(n2074), .Q(n1644) );
  MUX41X1 U2080 ( .IN1(reg5[8]), .IN3(reg7[8]), .IN2(reg6[8]), .IN4(reg8[8]), 
        .S0(n2033), .S1(n2074), .Q(n1645) );
  MUX41X1 U2081 ( .IN1(n1646), .IN3(n1644), .IN2(n1645), .IN4(n1643), .S0(
        n2011), .S1(n2017), .Q(n1647) );
  MUX21X1 U2082 ( .IN1(n1647), .IN2(n1642), .S(n2007), .Q(rd_dataB[8]) );
  MUX41X1 U2083 ( .IN1(reg29[9]), .IN3(reg31[9]), .IN2(reg30[9]), .IN4(
        reg32[9]), .S0(n2033), .S1(n2074), .Q(n1648) );
  MUX41X1 U2084 ( .IN1(reg25[9]), .IN3(reg27[9]), .IN2(reg26[9]), .IN4(
        reg28[9]), .S0(n2034), .S1(n2074), .Q(n1649) );
  MUX41X1 U2085 ( .IN1(reg21[9]), .IN3(reg23[9]), .IN2(reg22[9]), .IN4(
        reg24[9]), .S0(n2034), .S1(n2074), .Q(n1650) );
  MUX41X1 U2086 ( .IN1(reg17[9]), .IN3(reg19[9]), .IN2(reg18[9]), .IN4(
        reg20[9]), .S0(n2034), .S1(n2074), .Q(n1651) );
  MUX41X1 U2087 ( .IN1(n1651), .IN3(n1649), .IN2(n1650), .IN4(n1648), .S0(
        n2011), .S1(n2017), .Q(n1652) );
  MUX41X1 U2088 ( .IN1(reg13[9]), .IN3(reg15[9]), .IN2(reg14[9]), .IN4(
        reg16[9]), .S0(n2034), .S1(n2074), .Q(n1653) );
  MUX41X1 U2089 ( .IN1(reg9[9]), .IN3(reg11[9]), .IN2(reg10[9]), .IN4(reg12[9]), .S0(n2034), .S1(n2074), .Q(n1654) );
  MUX41X1 U2090 ( .IN1(reg5[9]), .IN3(reg7[9]), .IN2(reg6[9]), .IN4(reg8[9]), 
        .S0(n2034), .S1(n2074), .Q(n1655) );
  MUX41X1 U2091 ( .IN1(n1656), .IN3(n1654), .IN2(n1655), .IN4(n1653), .S0(
        n2011), .S1(n2017), .Q(n1657) );
  MUX21X1 U2092 ( .IN1(n1657), .IN2(n1652), .S(n2007), .Q(rd_dataB[9]) );
  MUX41X1 U2093 ( .IN1(reg29[10]), .IN3(reg31[10]), .IN2(reg30[10]), .IN4(
        reg32[10]), .S0(n2034), .S1(n2074), .Q(n1658) );
  MUX41X1 U2094 ( .IN1(reg25[10]), .IN3(reg27[10]), .IN2(reg26[10]), .IN4(
        reg28[10]), .S0(n2034), .S1(n2074), .Q(n1659) );
  MUX41X1 U2095 ( .IN1(reg21[10]), .IN3(reg23[10]), .IN2(reg22[10]), .IN4(
        reg24[10]), .S0(n2034), .S1(n2074), .Q(n1660) );
  MUX41X1 U2096 ( .IN1(reg17[10]), .IN3(reg19[10]), .IN2(reg18[10]), .IN4(
        reg20[10]), .S0(n2034), .S1(n2075), .Q(n1661) );
  MUX41X1 U2097 ( .IN1(n1661), .IN3(n1659), .IN2(n1660), .IN4(n1658), .S0(
        n2011), .S1(n2017), .Q(n1662) );
  MUX41X1 U2098 ( .IN1(reg13[10]), .IN3(reg15[10]), .IN2(reg14[10]), .IN4(
        reg16[10]), .S0(n2034), .S1(n2075), .Q(n1663) );
  MUX41X1 U2099 ( .IN1(reg9[10]), .IN3(reg11[10]), .IN2(reg10[10]), .IN4(
        reg12[10]), .S0(n2034), .S1(n2075), .Q(n1664) );
  MUX41X1 U2100 ( .IN1(reg5[10]), .IN3(reg7[10]), .IN2(reg6[10]), .IN4(
        reg8[10]), .S0(n2034), .S1(n2075), .Q(n1665) );
  MUX41X1 U2101 ( .IN1(n1666), .IN3(n1664), .IN2(n1665), .IN4(n1663), .S0(
        n2011), .S1(n2017), .Q(n1667) );
  MUX21X1 U2102 ( .IN1(n1667), .IN2(n1662), .S(n2007), .Q(rd_dataB[10]) );
  MUX41X1 U2103 ( .IN1(reg29[11]), .IN3(reg31[11]), .IN2(reg30[11]), .IN4(
        reg32[11]), .S0(n2034), .S1(n2075), .Q(n1668) );
  MUX41X1 U2104 ( .IN1(reg25[11]), .IN3(reg27[11]), .IN2(reg26[11]), .IN4(
        reg28[11]), .S0(n2035), .S1(n2075), .Q(n1669) );
  MUX41X1 U2105 ( .IN1(reg21[11]), .IN3(reg23[11]), .IN2(reg22[11]), .IN4(
        reg24[11]), .S0(n2035), .S1(n2075), .Q(n1670) );
  MUX41X1 U2106 ( .IN1(reg17[11]), .IN3(reg19[11]), .IN2(reg18[11]), .IN4(
        reg20[11]), .S0(n2035), .S1(n2075), .Q(n1671) );
  MUX41X1 U2107 ( .IN1(n1671), .IN3(n1669), .IN2(n1670), .IN4(n1668), .S0(
        n2011), .S1(n2017), .Q(n1672) );
  MUX41X1 U2108 ( .IN1(reg13[11]), .IN3(reg15[11]), .IN2(reg14[11]), .IN4(
        reg16[11]), .S0(n2035), .S1(n2075), .Q(n1673) );
  MUX41X1 U2109 ( .IN1(reg9[11]), .IN3(reg11[11]), .IN2(reg10[11]), .IN4(
        reg12[11]), .S0(n2035), .S1(n2075), .Q(n1674) );
  MUX41X1 U2110 ( .IN1(reg5[11]), .IN3(reg7[11]), .IN2(reg6[11]), .IN4(
        reg8[11]), .S0(n2035), .S1(n2075), .Q(n1675) );
  MUX41X1 U2111 ( .IN1(n1676), .IN3(n1674), .IN2(n1675), .IN4(n1673), .S0(
        n2011), .S1(n2017), .Q(n1677) );
  MUX21X1 U2112 ( .IN1(n1677), .IN2(n1672), .S(n2007), .Q(rd_dataB[11]) );
  MUX41X1 U2113 ( .IN1(reg29[12]), .IN3(reg31[12]), .IN2(reg30[12]), .IN4(
        reg32[12]), .S0(n2035), .S1(n2076), .Q(n1678) );
  MUX41X1 U2114 ( .IN1(reg25[12]), .IN3(reg27[12]), .IN2(reg26[12]), .IN4(
        reg28[12]), .S0(n2035), .S1(n2076), .Q(n1679) );
  MUX41X1 U2115 ( .IN1(reg21[12]), .IN3(reg23[12]), .IN2(reg22[12]), .IN4(
        reg24[12]), .S0(n2035), .S1(n2076), .Q(n1680) );
  MUX41X1 U2116 ( .IN1(reg17[12]), .IN3(reg19[12]), .IN2(reg18[12]), .IN4(
        reg20[12]), .S0(n2035), .S1(n2076), .Q(n1681) );
  MUX41X1 U2117 ( .IN1(n1681), .IN3(n1679), .IN2(n1680), .IN4(n1678), .S0(
        n2011), .S1(n2017), .Q(n1682) );
  MUX41X1 U2118 ( .IN1(reg13[12]), .IN3(reg15[12]), .IN2(reg14[12]), .IN4(
        reg16[12]), .S0(n2035), .S1(n2076), .Q(n1683) );
  MUX41X1 U2119 ( .IN1(reg9[12]), .IN3(reg11[12]), .IN2(reg10[12]), .IN4(
        reg12[12]), .S0(n2035), .S1(n2076), .Q(n1684) );
  MUX41X1 U2120 ( .IN1(reg5[12]), .IN3(reg7[12]), .IN2(reg6[12]), .IN4(
        reg8[12]), .S0(n2035), .S1(n2076), .Q(n1685) );
  MUX41X1 U2121 ( .IN1(n1686), .IN3(n1684), .IN2(n1685), .IN4(n1683), .S0(
        n2011), .S1(n2017), .Q(n1687) );
  MUX21X1 U2122 ( .IN1(n1687), .IN2(n1682), .S(n2007), .Q(rd_dataB[12]) );
  MUX41X1 U2123 ( .IN1(reg29[13]), .IN3(reg31[13]), .IN2(reg30[13]), .IN4(
        reg32[13]), .S0(n2035), .S1(n2076), .Q(n1688) );
  MUX41X1 U2124 ( .IN1(reg25[13]), .IN3(reg27[13]), .IN2(reg26[13]), .IN4(
        reg28[13]), .S0(n2035), .S1(n2076), .Q(n1689) );
  MUX41X1 U2125 ( .IN1(reg21[13]), .IN3(reg23[13]), .IN2(reg22[13]), .IN4(
        reg24[13]), .S0(n2036), .S1(n2076), .Q(n1690) );
  MUX41X1 U2126 ( .IN1(reg17[13]), .IN3(reg19[13]), .IN2(reg18[13]), .IN4(
        reg20[13]), .S0(n2036), .S1(n2076), .Q(n1691) );
  MUX41X1 U2127 ( .IN1(n1691), .IN3(n1689), .IN2(n1690), .IN4(n1688), .S0(
        n2011), .S1(n2017), .Q(n1692) );
  MUX41X1 U2128 ( .IN1(reg13[13]), .IN3(reg15[13]), .IN2(reg14[13]), .IN4(
        reg16[13]), .S0(n2036), .S1(n2076), .Q(n1693) );
  MUX41X1 U2129 ( .IN1(reg9[13]), .IN3(reg11[13]), .IN2(reg10[13]), .IN4(
        reg12[13]), .S0(n2036), .S1(n2077), .Q(n1694) );
  MUX41X1 U2130 ( .IN1(reg5[13]), .IN3(reg7[13]), .IN2(reg6[13]), .IN4(
        reg8[13]), .S0(n2036), .S1(n2078), .Q(n1695) );
  MUX41X1 U2131 ( .IN1(n1696), .IN3(n1694), .IN2(n1695), .IN4(n1693), .S0(
        n2011), .S1(n2017), .Q(n1697) );
  MUX21X1 U2132 ( .IN1(n1697), .IN2(n1692), .S(n2007), .Q(rd_dataB[13]) );
  MUX41X1 U2133 ( .IN1(reg29[14]), .IN3(reg31[14]), .IN2(reg30[14]), .IN4(
        reg32[14]), .S0(n2036), .S1(n2064), .Q(n1698) );
  MUX41X1 U2134 ( .IN1(reg25[14]), .IN3(reg27[14]), .IN2(reg26[14]), .IN4(
        reg28[14]), .S0(n2036), .S1(n2065), .Q(n1699) );
  MUX41X1 U2135 ( .IN1(reg21[14]), .IN3(reg23[14]), .IN2(reg22[14]), .IN4(
        reg24[14]), .S0(n2036), .S1(n2067), .Q(n1700) );
  MUX41X1 U2136 ( .IN1(reg17[14]), .IN3(reg19[14]), .IN2(reg18[14]), .IN4(
        reg20[14]), .S0(n2036), .S1(n2063), .Q(n1701) );
  MUX41X1 U2137 ( .IN1(n1701), .IN3(n1699), .IN2(n1700), .IN4(n1698), .S0(
        n2012), .S1(n2018), .Q(n1702) );
  MUX41X1 U2138 ( .IN1(reg13[14]), .IN3(reg15[14]), .IN2(reg14[14]), .IN4(
        reg16[14]), .S0(n2036), .S1(n2068), .Q(n1703) );
  MUX41X1 U2139 ( .IN1(reg9[14]), .IN3(reg11[14]), .IN2(reg10[14]), .IN4(
        reg12[14]), .S0(n2036), .S1(n2066), .Q(n1704) );
  MUX41X1 U2140 ( .IN1(reg5[14]), .IN3(reg7[14]), .IN2(reg6[14]), .IN4(
        reg8[14]), .S0(n2036), .S1(n2060), .Q(n1705) );
  MUX41X1 U2141 ( .IN1(n1706), .IN3(n1704), .IN2(n1705), .IN4(n1703), .S0(
        n2012), .S1(n2018), .Q(n1707) );
  MUX21X1 U2142 ( .IN1(n1707), .IN2(n1702), .S(n2007), .Q(rd_dataB[14]) );
  MUX41X1 U2143 ( .IN1(reg29[15]), .IN3(reg31[15]), .IN2(reg30[15]), .IN4(
        reg32[15]), .S0(n2037), .S1(n2067), .Q(n1708) );
  MUX41X1 U2144 ( .IN1(reg25[15]), .IN3(reg27[15]), .IN2(reg26[15]), .IN4(
        reg28[15]), .S0(n2037), .S1(n2068), .Q(n1709) );
  MUX41X1 U2145 ( .IN1(reg21[15]), .IN3(reg23[15]), .IN2(reg22[15]), .IN4(
        reg24[15]), .S0(n2036), .S1(n2066), .Q(n1710) );
  MUX41X1 U2146 ( .IN1(reg17[15]), .IN3(reg19[15]), .IN2(reg18[15]), .IN4(
        reg20[15]), .S0(n2037), .S1(n2077), .Q(n1711) );
  MUX41X1 U2147 ( .IN1(n1711), .IN3(n1709), .IN2(n1710), .IN4(n1708), .S0(
        n2012), .S1(n2018), .Q(n1712) );
  MUX41X1 U2148 ( .IN1(reg13[15]), .IN3(reg15[15]), .IN2(reg14[15]), .IN4(
        reg16[15]), .S0(n2037), .S1(n2077), .Q(n1713) );
  MUX41X1 U2149 ( .IN1(reg9[15]), .IN3(reg11[15]), .IN2(reg10[15]), .IN4(
        reg12[15]), .S0(n2036), .S1(n2077), .Q(n1714) );
  MUX41X1 U2150 ( .IN1(reg5[15]), .IN3(reg7[15]), .IN2(reg6[15]), .IN4(
        reg8[15]), .S0(n2037), .S1(n2077), .Q(n1715) );
  MUX41X1 U2151 ( .IN1(n1716), .IN3(n1714), .IN2(n1715), .IN4(n1713), .S0(
        n2012), .S1(n2018), .Q(n1717) );
  MUX21X1 U2152 ( .IN1(n1717), .IN2(n1712), .S(n2007), .Q(rd_dataB[15]) );
  MUX41X1 U2153 ( .IN1(reg29[16]), .IN3(reg31[16]), .IN2(reg30[16]), .IN4(
        reg32[16]), .S0(n2037), .S1(n2077), .Q(n1718) );
  MUX41X1 U2154 ( .IN1(reg25[16]), .IN3(reg27[16]), .IN2(reg26[16]), .IN4(
        reg28[16]), .S0(n2037), .S1(n2077), .Q(n1719) );
  MUX41X1 U2155 ( .IN1(reg21[16]), .IN3(reg23[16]), .IN2(reg22[16]), .IN4(
        reg24[16]), .S0(n2037), .S1(n2077), .Q(n1720) );
  MUX41X1 U2156 ( .IN1(reg17[16]), .IN3(reg19[16]), .IN2(reg18[16]), .IN4(
        reg20[16]), .S0(n2037), .S1(n2077), .Q(n1721) );
  MUX41X1 U2157 ( .IN1(n1721), .IN3(n1719), .IN2(n1720), .IN4(n1718), .S0(
        n2012), .S1(n2018), .Q(n1722) );
  MUX41X1 U2158 ( .IN1(reg13[16]), .IN3(reg15[16]), .IN2(reg14[16]), .IN4(
        reg16[16]), .S0(n2037), .S1(n2077), .Q(n1723) );
  MUX41X1 U2159 ( .IN1(reg9[16]), .IN3(reg11[16]), .IN2(reg10[16]), .IN4(
        reg12[16]), .S0(n2037), .S1(n2077), .Q(n1724) );
  MUX41X1 U2160 ( .IN1(reg5[16]), .IN3(reg7[16]), .IN2(reg6[16]), .IN4(
        reg8[16]), .S0(n2036), .S1(n2077), .Q(n1725) );
  MUX41X1 U2161 ( .IN1(n1726), .IN3(n1724), .IN2(n1725), .IN4(n1723), .S0(
        n2012), .S1(n2018), .Q(n1727) );
  MUX21X1 U2162 ( .IN1(n1727), .IN2(n1722), .S(n2007), .Q(rd_dataB[16]) );
  MUX41X1 U2163 ( .IN1(reg29[17]), .IN3(reg31[17]), .IN2(reg30[17]), .IN4(
        reg32[17]), .S0(n2037), .S1(n2077), .Q(n1728) );
  MUX41X1 U2164 ( .IN1(reg25[17]), .IN3(reg27[17]), .IN2(reg26[17]), .IN4(
        reg28[17]), .S0(n2037), .S1(n2078), .Q(n1729) );
  MUX41X1 U2165 ( .IN1(reg21[17]), .IN3(reg23[17]), .IN2(reg22[17]), .IN4(
        reg24[17]), .S0(n2038), .S1(n2078), .Q(n1730) );
  MUX41X1 U2166 ( .IN1(reg17[17]), .IN3(reg19[17]), .IN2(reg18[17]), .IN4(
        reg20[17]), .S0(n2037), .S1(n2078), .Q(n1731) );
  MUX41X1 U2167 ( .IN1(n1731), .IN3(n1729), .IN2(n1730), .IN4(n1728), .S0(
        n2012), .S1(n2018), .Q(n1732) );
  MUX41X1 U2168 ( .IN1(reg13[17]), .IN3(reg15[17]), .IN2(reg14[17]), .IN4(
        reg16[17]), .S0(n2038), .S1(n2078), .Q(n1733) );
  MUX41X1 U2169 ( .IN1(reg9[17]), .IN3(reg11[17]), .IN2(reg10[17]), .IN4(
        reg12[17]), .S0(n2038), .S1(n2078), .Q(n1734) );
  MUX41X1 U2170 ( .IN1(reg5[17]), .IN3(reg7[17]), .IN2(reg6[17]), .IN4(
        reg8[17]), .S0(n2037), .S1(n2078), .Q(n1735) );
  MUX41X1 U2171 ( .IN1(n1736), .IN3(n1734), .IN2(n1735), .IN4(n1733), .S0(
        n2012), .S1(n2018), .Q(n1737) );
  MUX21X1 U2172 ( .IN1(n1737), .IN2(n1732), .S(n2007), .Q(rd_dataB[17]) );
  MUX41X1 U2173 ( .IN1(reg29[18]), .IN3(reg31[18]), .IN2(reg30[18]), .IN4(
        reg32[18]), .S0(n2038), .S1(n2078), .Q(n1738) );
  MUX41X1 U2174 ( .IN1(reg25[18]), .IN3(reg27[18]), .IN2(reg26[18]), .IN4(
        reg28[18]), .S0(n2034), .S1(n2078), .Q(n1739) );
  MUX41X1 U2175 ( .IN1(reg21[18]), .IN3(reg23[18]), .IN2(reg22[18]), .IN4(
        reg24[18]), .S0(n2023), .S1(n2078), .Q(n1740) );
  MUX41X1 U2176 ( .IN1(reg17[18]), .IN3(reg19[18]), .IN2(reg18[18]), .IN4(
        reg20[18]), .S0(n2023), .S1(n2078), .Q(n1741) );
  MUX41X1 U2177 ( .IN1(n1741), .IN3(n1739), .IN2(n1740), .IN4(n1738), .S0(
        n2012), .S1(n2018), .Q(n1742) );
  MUX41X1 U2178 ( .IN1(reg13[18]), .IN3(reg15[18]), .IN2(reg14[18]), .IN4(
        reg16[18]), .S0(n2023), .S1(n2078), .Q(n1743) );
  MUX41X1 U2179 ( .IN1(reg9[18]), .IN3(reg11[18]), .IN2(reg10[18]), .IN4(
        reg12[18]), .S0(n2023), .S1(n2078), .Q(n1744) );
  MUX41X1 U2180 ( .IN1(reg5[18]), .IN3(reg7[18]), .IN2(reg6[18]), .IN4(
        reg8[18]), .S0(n2023), .S1(n2079), .Q(n1745) );
  MUX41X1 U2181 ( .IN1(n1746), .IN3(n1744), .IN2(n1745), .IN4(n1743), .S0(
        n2012), .S1(n2018), .Q(n1747) );
  MUX21X1 U2182 ( .IN1(n1747), .IN2(n1742), .S(n2007), .Q(rd_dataB[18]) );
  MUX41X1 U2183 ( .IN1(reg29[19]), .IN3(reg31[19]), .IN2(reg30[19]), .IN4(
        reg32[19]), .S0(n2023), .S1(n2079), .Q(n1748) );
  MUX41X1 U2184 ( .IN1(reg25[19]), .IN3(reg27[19]), .IN2(reg26[19]), .IN4(
        reg28[19]), .S0(n2023), .S1(n2079), .Q(n1749) );
  MUX41X1 U2185 ( .IN1(reg21[19]), .IN3(reg23[19]), .IN2(reg22[19]), .IN4(
        reg24[19]), .S0(n2023), .S1(n2079), .Q(n1750) );
  MUX41X1 U2186 ( .IN1(reg17[19]), .IN3(reg19[19]), .IN2(reg18[19]), .IN4(
        reg20[19]), .S0(n2023), .S1(n2079), .Q(n1751) );
  MUX41X1 U2187 ( .IN1(n1751), .IN3(n1749), .IN2(n1750), .IN4(n1748), .S0(
        n2012), .S1(n2018), .Q(n1752) );
  MUX41X1 U2188 ( .IN1(reg13[19]), .IN3(reg15[19]), .IN2(reg14[19]), .IN4(
        reg16[19]), .S0(n2024), .S1(n2079), .Q(n1753) );
  MUX41X1 U2189 ( .IN1(reg9[19]), .IN3(reg11[19]), .IN2(reg10[19]), .IN4(
        reg12[19]), .S0(n2024), .S1(n2079), .Q(n1754) );
  MUX41X1 U2190 ( .IN1(reg5[19]), .IN3(reg7[19]), .IN2(reg6[19]), .IN4(
        reg8[19]), .S0(n2024), .S1(n2079), .Q(n1755) );
  MUX41X1 U2191 ( .IN1(n1756), .IN3(n1754), .IN2(n1755), .IN4(n1753), .S0(
        n2012), .S1(n2018), .Q(n1757) );
  MUX21X1 U2192 ( .IN1(n1757), .IN2(n1752), .S(n2007), .Q(rd_dataB[19]) );
  MUX41X1 U2193 ( .IN1(reg29[20]), .IN3(reg31[20]), .IN2(reg30[20]), .IN4(
        reg32[20]), .S0(n2024), .S1(n2079), .Q(n1758) );
  MUX41X1 U2194 ( .IN1(reg25[20]), .IN3(reg27[20]), .IN2(reg26[20]), .IN4(
        reg28[20]), .S0(n2024), .S1(n2079), .Q(n1759) );
  MUX41X1 U2195 ( .IN1(reg21[20]), .IN3(reg23[20]), .IN2(reg22[20]), .IN4(
        reg24[20]), .S0(n2024), .S1(n2079), .Q(n1760) );
  MUX41X1 U2196 ( .IN1(reg17[20]), .IN3(reg19[20]), .IN2(reg18[20]), .IN4(
        reg20[20]), .S0(n2024), .S1(n2075), .Q(n1761) );
  MUX41X1 U2197 ( .IN1(n1761), .IN3(n1759), .IN2(n1760), .IN4(n1758), .S0(
        n2013), .S1(n2019), .Q(n1762) );
  MUX41X1 U2198 ( .IN1(reg13[20]), .IN3(reg15[20]), .IN2(reg14[20]), .IN4(
        reg16[20]), .S0(n2026), .S1(n2065), .Q(n1763) );
  MUX41X1 U2199 ( .IN1(reg9[20]), .IN3(reg11[20]), .IN2(reg10[20]), .IN4(
        reg12[20]), .S0(n2024), .S1(n2062), .Q(n1764) );
  MUX41X1 U2200 ( .IN1(reg5[20]), .IN3(reg7[20]), .IN2(reg6[20]), .IN4(
        reg8[20]), .S0(n2024), .S1(n2062), .Q(n1765) );
  MUX41X1 U2201 ( .IN1(n1766), .IN3(n1764), .IN2(n1765), .IN4(n1763), .S0(
        n2013), .S1(n2019), .Q(n1767) );
  MUX21X1 U2202 ( .IN1(n1767), .IN2(n1762), .S(n2008), .Q(rd_dataB[20]) );
  MUX41X1 U2203 ( .IN1(reg29[21]), .IN3(reg31[21]), .IN2(reg30[21]), .IN4(
        reg32[21]), .S0(n2024), .S1(n2062), .Q(n1768) );
  MUX41X1 U2204 ( .IN1(reg25[21]), .IN3(reg27[21]), .IN2(reg26[21]), .IN4(
        reg28[21]), .S0(n2024), .S1(n2062), .Q(n1769) );
  MUX41X1 U2205 ( .IN1(reg21[21]), .IN3(reg23[21]), .IN2(reg22[21]), .IN4(
        reg24[21]), .S0(n2024), .S1(n2062), .Q(n1770) );
  MUX41X1 U2206 ( .IN1(reg17[21]), .IN3(reg19[21]), .IN2(reg18[21]), .IN4(
        reg20[21]), .S0(n2024), .S1(n2062), .Q(n1771) );
  MUX41X1 U2207 ( .IN1(n1771), .IN3(n1769), .IN2(n1770), .IN4(n1768), .S0(
        n2013), .S1(n2019), .Q(n1772) );
  MUX41X1 U2208 ( .IN1(reg13[21]), .IN3(reg15[21]), .IN2(reg14[21]), .IN4(
        reg16[21]), .S0(n2024), .S1(n2062), .Q(n1773) );
  MUX41X1 U2209 ( .IN1(reg9[21]), .IN3(reg11[21]), .IN2(reg10[21]), .IN4(
        reg12[21]), .S0(n2025), .S1(n2063), .Q(n1774) );
  MUX41X1 U2210 ( .IN1(reg5[21]), .IN3(reg7[21]), .IN2(reg6[21]), .IN4(
        reg8[21]), .S0(n2025), .S1(n2063), .Q(n1775) );
  MUX41X1 U2211 ( .IN1(n1776), .IN3(n1774), .IN2(n1775), .IN4(n1773), .S0(
        n2013), .S1(n2019), .Q(n1777) );
  MUX21X1 U2212 ( .IN1(n1777), .IN2(n1772), .S(n2008), .Q(rd_dataB[21]) );
  MUX41X1 U2213 ( .IN1(reg29[22]), .IN3(reg31[22]), .IN2(reg30[22]), .IN4(
        reg32[22]), .S0(n2025), .S1(n2063), .Q(n1778) );
  MUX41X1 U2214 ( .IN1(reg25[22]), .IN3(reg27[22]), .IN2(reg26[22]), .IN4(
        reg28[22]), .S0(n2025), .S1(n2063), .Q(n1779) );
  MUX41X1 U2215 ( .IN1(reg21[22]), .IN3(reg23[22]), .IN2(reg22[22]), .IN4(
        reg24[22]), .S0(n2025), .S1(n2063), .Q(n1780) );
  MUX41X1 U2216 ( .IN1(reg17[22]), .IN3(reg19[22]), .IN2(reg18[22]), .IN4(
        reg20[22]), .S0(n2025), .S1(n2063), .Q(n1781) );
  MUX41X1 U2217 ( .IN1(n1781), .IN3(n1779), .IN2(n1780), .IN4(n1778), .S0(
        n2013), .S1(n2019), .Q(n1782) );
  MUX41X1 U2218 ( .IN1(reg13[22]), .IN3(reg15[22]), .IN2(reg14[22]), .IN4(
        reg16[22]), .S0(n2025), .S1(n2063), .Q(n1783) );
  MUX41X1 U2219 ( .IN1(reg9[22]), .IN3(reg11[22]), .IN2(reg10[22]), .IN4(
        reg12[22]), .S0(n2025), .S1(n2063), .Q(n1784) );
  MUX41X1 U2220 ( .IN1(reg5[22]), .IN3(reg7[22]), .IN2(reg6[22]), .IN4(
        reg8[22]), .S0(n2025), .S1(n2063), .Q(n1785) );
  MUX41X1 U2221 ( .IN1(n1786), .IN3(n1784), .IN2(n1785), .IN4(n1783), .S0(
        n2013), .S1(n2019), .Q(n1787) );
  MUX21X1 U2222 ( .IN1(n1787), .IN2(n1782), .S(n2008), .Q(rd_dataB[22]) );
  MUX41X1 U2223 ( .IN1(reg29[23]), .IN3(reg31[23]), .IN2(reg30[23]), .IN4(
        reg32[23]), .S0(n2025), .S1(n2063), .Q(n1788) );
  MUX41X1 U2224 ( .IN1(reg25[23]), .IN3(reg27[23]), .IN2(reg26[23]), .IN4(
        reg28[23]), .S0(n2025), .S1(n2063), .Q(n1789) );
  MUX41X1 U2225 ( .IN1(reg21[23]), .IN3(reg23[23]), .IN2(reg22[23]), .IN4(
        reg24[23]), .S0(n2025), .S1(n2063), .Q(n1790) );
  MUX41X1 U2226 ( .IN1(reg17[23]), .IN3(reg19[23]), .IN2(reg18[23]), .IN4(
        reg20[23]), .S0(n2025), .S1(n2064), .Q(n1791) );
  MUX41X1 U2227 ( .IN1(n1791), .IN3(n1789), .IN2(n1790), .IN4(n1788), .S0(
        n2013), .S1(n2019), .Q(n1792) );
  MUX41X1 U2228 ( .IN1(reg13[23]), .IN3(reg15[23]), .IN2(reg14[23]), .IN4(
        reg16[23]), .S0(n2025), .S1(n2064), .Q(n1793) );
  MUX41X1 U2229 ( .IN1(reg9[23]), .IN3(reg11[23]), .IN2(reg10[23]), .IN4(
        reg12[23]), .S0(n2025), .S1(n2064), .Q(n1794) );
  MUX41X1 U2230 ( .IN1(reg5[23]), .IN3(reg7[23]), .IN2(reg6[23]), .IN4(
        reg8[23]), .S0(n2026), .S1(n2064), .Q(n1795) );
  MUX41X1 U2231 ( .IN1(n1796), .IN3(n1794), .IN2(n1795), .IN4(n1793), .S0(
        n2013), .S1(n2019), .Q(n1797) );
  MUX21X1 U2232 ( .IN1(n1797), .IN2(n1792), .S(n2008), .Q(rd_dataB[23]) );
  MUX41X1 U2233 ( .IN1(reg29[24]), .IN3(reg31[24]), .IN2(reg30[24]), .IN4(
        reg32[24]), .S0(n2026), .S1(n2064), .Q(n1798) );
  MUX41X1 U2234 ( .IN1(reg25[24]), .IN3(reg27[24]), .IN2(reg26[24]), .IN4(
        reg28[24]), .S0(n2026), .S1(n2064), .Q(n1799) );
  MUX41X1 U2235 ( .IN1(reg21[24]), .IN3(reg23[24]), .IN2(reg22[24]), .IN4(
        reg24[24]), .S0(n2026), .S1(n2064), .Q(n1800) );
  MUX41X1 U2236 ( .IN1(reg17[24]), .IN3(reg19[24]), .IN2(reg18[24]), .IN4(
        reg20[24]), .S0(n2026), .S1(n2064), .Q(n1801) );
  MUX41X1 U2237 ( .IN1(n1801), .IN3(n1799), .IN2(n1800), .IN4(n1798), .S0(
        n2013), .S1(n2019), .Q(n1802) );
  MUX41X1 U2238 ( .IN1(reg13[24]), .IN3(reg15[24]), .IN2(reg14[24]), .IN4(
        reg16[24]), .S0(n2026), .S1(n2064), .Q(n1803) );
  MUX41X1 U2239 ( .IN1(reg9[24]), .IN3(reg11[24]), .IN2(reg10[24]), .IN4(
        reg12[24]), .S0(n2026), .S1(n2064), .Q(n1804) );
  MUX41X1 U2240 ( .IN1(reg5[24]), .IN3(reg7[24]), .IN2(reg6[24]), .IN4(
        reg8[24]), .S0(n2026), .S1(n2064), .Q(n1805) );
  MUX41X1 U2241 ( .IN1(n1806), .IN3(n1804), .IN2(n1805), .IN4(n1803), .S0(
        n2013), .S1(n2019), .Q(n1807) );
  MUX21X1 U2242 ( .IN1(n1807), .IN2(n1802), .S(n2008), .Q(rd_dataB[24]) );
  MUX41X1 U2243 ( .IN1(reg29[25]), .IN3(reg31[25]), .IN2(reg30[25]), .IN4(
        reg32[25]), .S0(n2026), .S1(n2064), .Q(n1808) );
  MUX41X1 U2244 ( .IN1(reg25[25]), .IN3(reg27[25]), .IN2(reg26[25]), .IN4(
        reg28[25]), .S0(n2026), .S1(n2065), .Q(n1809) );
  MUX41X1 U2245 ( .IN1(reg21[25]), .IN3(reg23[25]), .IN2(reg22[25]), .IN4(
        reg24[25]), .S0(n2026), .S1(n2065), .Q(n1810) );
  MUX41X1 U2246 ( .IN1(reg17[25]), .IN3(reg19[25]), .IN2(reg18[25]), .IN4(
        reg20[25]), .S0(n2026), .S1(n2065), .Q(n1811) );
  MUX41X1 U2247 ( .IN1(n1811), .IN3(n1809), .IN2(n1810), .IN4(n1808), .S0(
        n2013), .S1(n2019), .Q(n1812) );
  MUX41X1 U2248 ( .IN1(reg13[25]), .IN3(reg15[25]), .IN2(reg14[25]), .IN4(
        reg16[25]), .S0(n2026), .S1(n2065), .Q(n1813) );
  MUX41X1 U2249 ( .IN1(reg9[25]), .IN3(reg11[25]), .IN2(reg10[25]), .IN4(
        reg12[25]), .S0(n2026), .S1(n2065), .Q(n1814) );
  MUX41X1 U2250 ( .IN1(reg5[25]), .IN3(reg7[25]), .IN2(reg6[25]), .IN4(
        reg8[25]), .S0(n2027), .S1(n2065), .Q(n1815) );
  MUX41X1 U2251 ( .IN1(n1816), .IN3(n1814), .IN2(n1815), .IN4(n1813), .S0(
        n2013), .S1(n2019), .Q(n1817) );
  MUX21X1 U2252 ( .IN1(n1817), .IN2(n1812), .S(n2008), .Q(rd_dataB[25]) );
  MUX41X1 U2253 ( .IN1(reg29[26]), .IN3(reg31[26]), .IN2(reg30[26]), .IN4(
        reg32[26]), .S0(n2027), .S1(n2065), .Q(n1818) );
  MUX41X1 U2254 ( .IN1(reg25[26]), .IN3(reg27[26]), .IN2(reg26[26]), .IN4(
        reg28[26]), .S0(n2027), .S1(n2065), .Q(n1819) );
  MUX41X1 U2255 ( .IN1(reg21[26]), .IN3(reg23[26]), .IN2(reg22[26]), .IN4(
        reg24[26]), .S0(n2027), .S1(n2065), .Q(n1820) );
  MUX41X1 U2256 ( .IN1(reg17[26]), .IN3(reg19[26]), .IN2(reg18[26]), .IN4(
        reg20[26]), .S0(n2027), .S1(n2065), .Q(n1821) );
  MUX41X1 U2257 ( .IN1(n1821), .IN3(n1819), .IN2(n1820), .IN4(n1818), .S0(
        n2014), .S1(n2020), .Q(n1822) );
  MUX41X1 U2258 ( .IN1(reg13[26]), .IN3(reg15[26]), .IN2(reg14[26]), .IN4(
        reg16[26]), .S0(n2027), .S1(n2065), .Q(n1823) );
  MUX41X1 U2259 ( .IN1(reg9[26]), .IN3(reg11[26]), .IN2(reg10[26]), .IN4(
        reg12[26]), .S0(n2027), .S1(n2066), .Q(n1824) );
  MUX41X1 U2260 ( .IN1(reg5[26]), .IN3(reg7[26]), .IN2(reg6[26]), .IN4(
        reg8[26]), .S0(n2027), .S1(n2066), .Q(n1825) );
  MUX41X1 U2261 ( .IN1(n1826), .IN3(n1824), .IN2(n1825), .IN4(n1823), .S0(
        n2014), .S1(n2020), .Q(n1827) );
  MUX21X1 U2262 ( .IN1(n1827), .IN2(n1822), .S(n2008), .Q(rd_dataB[26]) );
  MUX41X1 U2263 ( .IN1(reg29[27]), .IN3(reg31[27]), .IN2(reg30[27]), .IN4(
        reg32[27]), .S0(n2027), .S1(n2066), .Q(n1828) );
  MUX41X1 U2264 ( .IN1(reg25[27]), .IN3(reg27[27]), .IN2(reg26[27]), .IN4(
        reg28[27]), .S0(n2027), .S1(n2066), .Q(n1829) );
  MUX41X1 U2265 ( .IN1(reg21[27]), .IN3(reg23[27]), .IN2(reg22[27]), .IN4(
        reg24[27]), .S0(n2027), .S1(n2066), .Q(n1830) );
  MUX41X1 U2266 ( .IN1(reg17[27]), .IN3(reg19[27]), .IN2(reg18[27]), .IN4(
        reg20[27]), .S0(n2027), .S1(n2066), .Q(n1831) );
  MUX41X1 U2267 ( .IN1(n1831), .IN3(n1829), .IN2(n1830), .IN4(n1828), .S0(
        n2014), .S1(n2020), .Q(n1832) );
  MUX41X1 U2268 ( .IN1(reg13[27]), .IN3(reg15[27]), .IN2(reg14[27]), .IN4(
        reg16[27]), .S0(n2027), .S1(n2066), .Q(n1833) );
  MUX41X1 U2269 ( .IN1(reg9[27]), .IN3(reg11[27]), .IN2(reg10[27]), .IN4(
        reg12[27]), .S0(n2027), .S1(n2066), .Q(n1834) );
  MUX41X1 U2270 ( .IN1(reg5[27]), .IN3(reg7[27]), .IN2(reg6[27]), .IN4(
        reg8[27]), .S0(n2027), .S1(n2066), .Q(n1835) );
  MUX41X1 U2271 ( .IN1(n1836), .IN3(n1834), .IN2(n1835), .IN4(n1833), .S0(
        n2014), .S1(n2020), .Q(n1837) );
  MUX21X1 U2272 ( .IN1(n1837), .IN2(n1832), .S(n2008), .Q(rd_dataB[27]) );
  MUX41X1 U2273 ( .IN1(reg29[28]), .IN3(reg31[28]), .IN2(reg30[28]), .IN4(
        reg32[28]), .S0(n2028), .S1(n2066), .Q(n1838) );
  MUX41X1 U2274 ( .IN1(reg25[28]), .IN3(reg27[28]), .IN2(reg26[28]), .IN4(
        reg28[28]), .S0(n2028), .S1(n2066), .Q(n1839) );
  MUX41X1 U2275 ( .IN1(reg21[28]), .IN3(reg23[28]), .IN2(reg22[28]), .IN4(
        reg24[28]), .S0(n2028), .S1(n2066), .Q(n1840) );
  MUX41X1 U2276 ( .IN1(reg17[28]), .IN3(reg19[28]), .IN2(reg18[28]), .IN4(
        reg20[28]), .S0(n2028), .S1(n2067), .Q(n1841) );
  MUX41X1 U2277 ( .IN1(n1841), .IN3(n1839), .IN2(n1840), .IN4(n1838), .S0(
        n2014), .S1(n2020), .Q(n1842) );
  MUX41X1 U2278 ( .IN1(reg13[28]), .IN3(reg15[28]), .IN2(reg14[28]), .IN4(
        reg16[28]), .S0(n2028), .S1(n2067), .Q(n1843) );
  MUX41X1 U2279 ( .IN1(reg9[28]), .IN3(reg11[28]), .IN2(reg10[28]), .IN4(
        reg12[28]), .S0(n2028), .S1(n2067), .Q(n1844) );
  MUX41X1 U2280 ( .IN1(reg5[28]), .IN3(reg7[28]), .IN2(reg6[28]), .IN4(
        reg8[28]), .S0(n2028), .S1(n2067), .Q(n1845) );
  MUX41X1 U2281 ( .IN1(n1846), .IN3(n1844), .IN2(n1845), .IN4(n1843), .S0(
        n2014), .S1(n2020), .Q(n1847) );
  MUX21X1 U2282 ( .IN1(n1847), .IN2(n1842), .S(n2008), .Q(rd_dataB[28]) );
  MUX41X1 U2283 ( .IN1(reg29[29]), .IN3(reg31[29]), .IN2(reg30[29]), .IN4(
        reg32[29]), .S0(n2028), .S1(n2067), .Q(n1848) );
  MUX41X1 U2284 ( .IN1(reg25[29]), .IN3(reg27[29]), .IN2(reg26[29]), .IN4(
        reg28[29]), .S0(n2028), .S1(n2067), .Q(n1849) );
  MUX41X1 U2285 ( .IN1(reg21[29]), .IN3(reg23[29]), .IN2(reg22[29]), .IN4(
        reg24[29]), .S0(n2028), .S1(n2067), .Q(n1850) );
  MUX41X1 U2286 ( .IN1(reg17[29]), .IN3(reg19[29]), .IN2(reg18[29]), .IN4(
        reg20[29]), .S0(n2028), .S1(n2067), .Q(n1851) );
  MUX41X1 U2287 ( .IN1(n1851), .IN3(n1849), .IN2(n1850), .IN4(n1848), .S0(
        n2014), .S1(n2020), .Q(n1852) );
  MUX41X1 U2288 ( .IN1(reg13[29]), .IN3(reg15[29]), .IN2(reg14[29]), .IN4(
        reg16[29]), .S0(n2028), .S1(n2067), .Q(n1853) );
  MUX41X1 U2289 ( .IN1(reg9[29]), .IN3(reg11[29]), .IN2(reg10[29]), .IN4(
        reg12[29]), .S0(n2028), .S1(n2067), .Q(n1854) );
  MUX41X1 U2290 ( .IN1(reg5[29]), .IN3(reg7[29]), .IN2(reg6[29]), .IN4(
        reg8[29]), .S0(n2028), .S1(n2067), .Q(n1855) );
  MUX41X1 U2291 ( .IN1(n1856), .IN3(n1854), .IN2(n1855), .IN4(n1853), .S0(
        n2014), .S1(n2020), .Q(n1857) );
  MUX21X1 U2292 ( .IN1(n1857), .IN2(n1852), .S(n2008), .Q(rd_dataB[29]) );
  MUX41X1 U2293 ( .IN1(reg29[30]), .IN3(reg31[30]), .IN2(reg30[30]), .IN4(
        reg32[30]), .S0(n2028), .S1(n2067), .Q(n1858) );
  MUX41X1 U2294 ( .IN1(reg25[30]), .IN3(reg27[30]), .IN2(reg26[30]), .IN4(
        reg28[30]), .S0(n2029), .S1(n2068), .Q(n1859) );
  MUX41X1 U2295 ( .IN1(reg21[30]), .IN3(reg23[30]), .IN2(reg22[30]), .IN4(
        reg24[30]), .S0(n2029), .S1(n2068), .Q(n1860) );
  MUX41X1 U2296 ( .IN1(reg17[30]), .IN3(reg19[30]), .IN2(reg18[30]), .IN4(
        reg20[30]), .S0(n2029), .S1(n2068), .Q(n1861) );
  MUX41X1 U2297 ( .IN1(n1861), .IN3(n1859), .IN2(n1860), .IN4(n1858), .S0(
        n2014), .S1(n2020), .Q(n1862) );
  MUX41X1 U2298 ( .IN1(reg13[30]), .IN3(reg15[30]), .IN2(reg14[30]), .IN4(
        reg16[30]), .S0(n2029), .S1(n2068), .Q(n1863) );
  MUX41X1 U2299 ( .IN1(reg9[30]), .IN3(reg11[30]), .IN2(reg10[30]), .IN4(
        reg12[30]), .S0(n2029), .S1(n2068), .Q(n1864) );
  MUX41X1 U2300 ( .IN1(reg5[30]), .IN3(reg7[30]), .IN2(reg6[30]), .IN4(
        reg8[30]), .S0(n2029), .S1(n2068), .Q(n1865) );
  MUX41X1 U2301 ( .IN1(n1866), .IN3(n1864), .IN2(n1865), .IN4(n1863), .S0(
        n2014), .S1(n2020), .Q(n1867) );
  MUX21X1 U2302 ( .IN1(n1867), .IN2(n1862), .S(n2008), .Q(rd_dataB[30]) );
  MUX41X1 U2303 ( .IN1(reg29[31]), .IN3(reg31[31]), .IN2(reg30[31]), .IN4(
        reg32[31]), .S0(n2029), .S1(n2068), .Q(n1868) );
  MUX41X1 U2304 ( .IN1(reg25[31]), .IN3(reg27[31]), .IN2(reg26[31]), .IN4(
        reg28[31]), .S0(n2029), .S1(n2068), .Q(n1869) );
  MUX41X1 U2305 ( .IN1(reg21[31]), .IN3(reg23[31]), .IN2(reg22[31]), .IN4(
        reg24[31]), .S0(n2029), .S1(n2068), .Q(n1870) );
  MUX41X1 U2306 ( .IN1(reg17[31]), .IN3(reg19[31]), .IN2(reg18[31]), .IN4(
        reg20[31]), .S0(n2029), .S1(n2068), .Q(n1871) );
  MUX41X1 U2307 ( .IN1(n1871), .IN3(n1869), .IN2(n1870), .IN4(n1868), .S0(
        n2014), .S1(n2020), .Q(n1872) );
  MUX41X1 U2308 ( .IN1(reg13[31]), .IN3(reg15[31]), .IN2(reg14[31]), .IN4(
        reg16[31]), .S0(n2029), .S1(n2068), .Q(n1873) );
  MUX41X1 U2309 ( .IN1(reg9[31]), .IN3(reg11[31]), .IN2(reg10[31]), .IN4(
        reg12[31]), .S0(n2029), .S1(n2068), .Q(n1874) );
  MUX41X1 U2310 ( .IN1(reg5[31]), .IN3(reg7[31]), .IN2(reg6[31]), .IN4(
        reg8[31]), .S0(n2029), .S1(n2069), .Q(n1875) );
  MUX41X1 U2311 ( .IN1(n1876), .IN3(n1874), .IN2(n1875), .IN4(n1873), .S0(
        n2014), .S1(n2020), .Q(n1877) );
  MUX21X1 U2312 ( .IN1(n1877), .IN2(n1872), .S(n2008), .Q(rd_dataB[31]) );
  MUX21X1 U2313 ( .IN1(n1878), .IN2(n1879), .S(n2038), .Q(n1881) );
  NAND3X0 U2314 ( .IN1(reg4[31]), .IN2(n2023), .IN3(n2058), .QN(n1880) );
  MUX21X1 U2315 ( .IN1(n1882), .IN2(n1883), .S(n2039), .Q(n1885) );
  NAND3X0 U2316 ( .IN1(reg4[30]), .IN2(n2023), .IN3(n2058), .QN(n1884) );
  MUX21X1 U2317 ( .IN1(n1886), .IN2(n1887), .S(n2038), .Q(n1889) );
  NAND3X0 U2318 ( .IN1(reg4[29]), .IN2(n2023), .IN3(n2058), .QN(n1888) );
  MUX21X1 U2319 ( .IN1(n1890), .IN2(n1891), .S(n2038), .Q(n1893) );
  NAND3X0 U2320 ( .IN1(reg4[28]), .IN2(n2023), .IN3(n2059), .QN(n1892) );
  MUX21X1 U2321 ( .IN1(n1894), .IN2(n1895), .S(n2039), .Q(n1897) );
  NAND3X0 U2322 ( .IN1(reg4[27]), .IN2(n2023), .IN3(n2059), .QN(n1896) );
  MUX21X1 U2323 ( .IN1(n1898), .IN2(n1899), .S(n2038), .Q(n1901) );
  NAND3X0 U2324 ( .IN1(reg4[26]), .IN2(n2023), .IN3(n2059), .QN(n1900) );
  MUX21X1 U2325 ( .IN1(n1902), .IN2(n1903), .S(n2038), .Q(n1905) );
  NAND3X0 U2326 ( .IN1(reg4[25]), .IN2(n2023), .IN3(n2059), .QN(n1904) );
  MUX21X1 U2327 ( .IN1(n1906), .IN2(n1907), .S(n2039), .Q(n1909) );
  NAND3X0 U2328 ( .IN1(reg4[24]), .IN2(n2022), .IN3(n2059), .QN(n1908) );
  MUX21X1 U2329 ( .IN1(n1910), .IN2(n1911), .S(n2038), .Q(n1913) );
  NAND3X0 U2330 ( .IN1(reg4[23]), .IN2(n2022), .IN3(n2059), .QN(n1912) );
  MUX21X1 U2331 ( .IN1(n1914), .IN2(n1915), .S(n2038), .Q(n1917) );
  NAND3X0 U2332 ( .IN1(reg4[22]), .IN2(n2022), .IN3(n2059), .QN(n1916) );
  MUX21X1 U2333 ( .IN1(n1918), .IN2(n1919), .S(n2039), .Q(n1921) );
  NAND3X0 U2334 ( .IN1(reg4[21]), .IN2(n2022), .IN3(n2059), .QN(n1920) );
  MUX21X1 U2335 ( .IN1(n1922), .IN2(n1923), .S(n2038), .Q(n1925) );
  NAND3X0 U2336 ( .IN1(reg4[20]), .IN2(n2022), .IN3(n2059), .QN(n1924) );
  MUX21X1 U2337 ( .IN1(n1926), .IN2(n1927), .S(n2039), .Q(n1929) );
  NAND3X0 U2338 ( .IN1(reg4[19]), .IN2(n2022), .IN3(n2059), .QN(n1928) );
  MUX21X1 U2339 ( .IN1(n1930), .IN2(n1931), .S(n2039), .Q(n1933) );
  NAND3X0 U2340 ( .IN1(reg4[18]), .IN2(n2022), .IN3(n2059), .QN(n1932) );
  MUX21X1 U2341 ( .IN1(n1934), .IN2(n1935), .S(n2039), .Q(n1937) );
  NAND3X0 U2342 ( .IN1(reg4[17]), .IN2(n2022), .IN3(n2059), .QN(n1936) );
  MUX21X1 U2343 ( .IN1(n1938), .IN2(n1939), .S(n2039), .Q(n1941) );
  NAND3X0 U2344 ( .IN1(reg4[16]), .IN2(n2022), .IN3(n2059), .QN(n1940) );
  MUX21X1 U2345 ( .IN1(n1942), .IN2(n1943), .S(n2040), .Q(n1945) );
  NAND3X0 U2346 ( .IN1(reg4[15]), .IN2(n2022), .IN3(n2059), .QN(n1944) );
  MUX21X1 U2347 ( .IN1(n1946), .IN2(n1947), .S(n2039), .Q(n1949) );
  NAND3X0 U2348 ( .IN1(reg4[14]), .IN2(n2022), .IN3(n2059), .QN(n1948) );
  MUX21X1 U2349 ( .IN1(n1950), .IN2(n1951), .S(n2039), .Q(n1953) );
  NAND3X0 U2350 ( .IN1(reg4[13]), .IN2(n2022), .IN3(n2059), .QN(n1952) );
  MUX21X1 U2351 ( .IN1(n1954), .IN2(n1955), .S(n2040), .Q(n1957) );
  NAND3X0 U2352 ( .IN1(reg4[12]), .IN2(n2022), .IN3(n2059), .QN(n1956) );
  MUX21X1 U2353 ( .IN1(n1958), .IN2(n1959), .S(n2039), .Q(n1961) );
  NAND3X0 U2354 ( .IN1(reg4[11]), .IN2(n2022), .IN3(n2059), .QN(n1960) );
  MUX21X1 U2355 ( .IN1(n1962), .IN2(n1963), .S(n2039), .Q(n1965) );
  NAND3X0 U2356 ( .IN1(reg4[10]), .IN2(n2022), .IN3(n2059), .QN(n1964) );
  MUX21X1 U2357 ( .IN1(n1966), .IN2(n1967), .S(n2040), .Q(n1969) );
  NAND3X0 U2358 ( .IN1(reg4[9]), .IN2(n2022), .IN3(n2059), .QN(n1968) );
  MUX21X1 U2359 ( .IN1(n1970), .IN2(n1971), .S(n2040), .Q(n1973) );
  NAND3X0 U2360 ( .IN1(reg4[8]), .IN2(n2022), .IN3(n2059), .QN(n1972) );
  MUX21X1 U2361 ( .IN1(n1974), .IN2(n1975), .S(n2040), .Q(n1977) );
  NAND3X0 U2362 ( .IN1(reg4[7]), .IN2(n2022), .IN3(n2059), .QN(n1976) );
  MUX21X1 U2363 ( .IN1(n1978), .IN2(n1979), .S(n2040), .Q(n1981) );
  NAND3X0 U2364 ( .IN1(reg4[6]), .IN2(n2021), .IN3(n2058), .QN(n1980) );
  MUX21X1 U2365 ( .IN1(n1982), .IN2(n1983), .S(n2040), .Q(n1985) );
  NAND3X0 U2366 ( .IN1(reg4[5]), .IN2(n2021), .IN3(n2059), .QN(n1984) );
  MUX21X1 U2367 ( .IN1(n1986), .IN2(n1987), .S(n2040), .Q(n1989) );
  NAND3X0 U2368 ( .IN1(reg4[4]), .IN2(n2021), .IN3(n2058), .QN(n1988) );
  MUX21X1 U2369 ( .IN1(n1990), .IN2(n1991), .S(n2040), .Q(n1993) );
  NAND3X0 U2370 ( .IN1(reg4[3]), .IN2(n2021), .IN3(n2058), .QN(n1992) );
  MUX21X1 U2371 ( .IN1(n1994), .IN2(n1995), .S(n2040), .Q(n1997) );
  NAND3X0 U2372 ( .IN1(reg4[2]), .IN2(n2021), .IN3(n2058), .QN(n1996) );
  MUX21X1 U2373 ( .IN1(n1998), .IN2(n1999), .S(n2040), .Q(n2001) );
  NAND3X0 U2374 ( .IN1(reg4[1]), .IN2(n2021), .IN3(n2058), .QN(n2000) );
  MUX21X1 U2375 ( .IN1(n2002), .IN2(n2003), .S(n2040), .Q(n2005) );
  NAND3X0 U2376 ( .IN1(reg4[0]), .IN2(n2021), .IN3(n2059), .QN(n2004) );
  INVX0 U2377 ( .INP(N16), .ZN(n2043) );
  INVX0 U2378 ( .INP(n2044), .ZN(n2058) );
  INVX0 U2379 ( .INP(n2045), .ZN(n2060) );
  INVX0 U2380 ( .INP(n2045), .ZN(n2061) );
  INVX0 U2381 ( .INP(n2045), .ZN(n2062) );
  INVX0 U2382 ( .INP(n2045), .ZN(n2063) );
  INVX0 U2383 ( .INP(n2045), .ZN(n2064) );
  INVX0 U2384 ( .INP(n2045), .ZN(n2065) );
  INVX0 U2385 ( .INP(n2045), .ZN(n2066) );
  INVX0 U2386 ( .INP(n2045), .ZN(n2067) );
  INVX0 U2387 ( .INP(n2045), .ZN(n2068) );
  INVX0 U2388 ( .INP(n2046), .ZN(n2069) );
  INVX0 U2389 ( .INP(n2046), .ZN(n2070) );
  INVX0 U2390 ( .INP(n2046), .ZN(n2071) );
  INVX0 U2391 ( .INP(n2046), .ZN(n2072) );
  INVX0 U2392 ( .INP(n2046), .ZN(n2073) );
  INVX0 U2393 ( .INP(n2046), .ZN(n2074) );
  INVX0 U2394 ( .INP(n2046), .ZN(n2075) );
  INVX0 U2395 ( .INP(n2046), .ZN(n2076) );
  NBUFFX4 U2396 ( .INP(n2043), .Z(n2045) );
  INVX0 U2397 ( .INP(n2082), .ZN(n2080) );
  INVX0 U2398 ( .INP(n2083), .ZN(n2081) );
  INVX0 U2399 ( .INP(n2086), .ZN(n2084) );
  INVX0 U2400 ( .INP(n2087), .ZN(n2085) );
  INVX0 U2401 ( .INP(n2090), .ZN(n2088) );
  INVX0 U2402 ( .INP(n2091), .ZN(n2089) );
  INVX0 U2403 ( .INP(n2094), .ZN(n2092) );
  INVX0 U2404 ( .INP(n2095), .ZN(n2093) );
  INVX0 U2405 ( .INP(n2098), .ZN(n2096) );
  INVX0 U2406 ( .INP(n2099), .ZN(n2097) );
  INVX0 U2407 ( .INP(n2102), .ZN(n2100) );
  INVX0 U2408 ( .INP(n2103), .ZN(n2101) );
  INVX0 U2409 ( .INP(n2106), .ZN(n2104) );
  INVX0 U2410 ( .INP(n2107), .ZN(n2105) );
  INVX0 U2411 ( .INP(n2110), .ZN(n2108) );
  INVX0 U2412 ( .INP(n2111), .ZN(n2109) );
  INVX0 U2413 ( .INP(n2114), .ZN(n2112) );
  INVX0 U2414 ( .INP(n2115), .ZN(n2113) );
  INVX0 U2415 ( .INP(n2118), .ZN(n2116) );
  INVX0 U2416 ( .INP(n2119), .ZN(n2117) );
  INVX0 U2417 ( .INP(n2122), .ZN(n2120) );
  INVX0 U2418 ( .INP(n2123), .ZN(n2121) );
  INVX0 U2419 ( .INP(n2126), .ZN(n2124) );
  INVX0 U2420 ( .INP(n2127), .ZN(n2125) );
  INVX0 U2421 ( .INP(n2130), .ZN(n2128) );
  INVX0 U2422 ( .INP(n2131), .ZN(n2129) );
  INVX0 U2423 ( .INP(n2134), .ZN(n2132) );
  INVX0 U2424 ( .INP(n2135), .ZN(n2133) );
  INVX0 U2425 ( .INP(n2138), .ZN(n2136) );
  INVX0 U2426 ( .INP(n2139), .ZN(n2137) );
  INVX0 U2427 ( .INP(n2142), .ZN(n2140) );
  INVX0 U2428 ( .INP(n2143), .ZN(n2141) );
  INVX0 U2429 ( .INP(n2146), .ZN(n2144) );
  INVX0 U2430 ( .INP(n2147), .ZN(n2145) );
  INVX0 U2431 ( .INP(n2150), .ZN(n2148) );
  INVX0 U2432 ( .INP(n2151), .ZN(n2149) );
  INVX0 U2433 ( .INP(n2154), .ZN(n2152) );
  INVX0 U2434 ( .INP(n2155), .ZN(n2153) );
  INVX0 U2435 ( .INP(n2158), .ZN(n2156) );
  INVX0 U2436 ( .INP(n2159), .ZN(n2157) );
  INVX0 U2437 ( .INP(n2162), .ZN(n2160) );
  INVX0 U2438 ( .INP(n2163), .ZN(n2161) );
  INVX0 U2439 ( .INP(n2166), .ZN(n2164) );
  INVX0 U2440 ( .INP(n2167), .ZN(n2165) );
  INVX0 U2441 ( .INP(n2170), .ZN(n2168) );
  INVX0 U2442 ( .INP(n2171), .ZN(n2169) );
  INVX0 U2443 ( .INP(n2174), .ZN(n2172) );
  INVX0 U2444 ( .INP(n2175), .ZN(n2173) );
  INVX0 U2445 ( .INP(n2178), .ZN(n2176) );
  INVX0 U2446 ( .INP(n2179), .ZN(n2177) );
  INVX0 U2447 ( .INP(n2182), .ZN(n2180) );
  INVX0 U2448 ( .INP(n2183), .ZN(n2181) );
  INVX0 U2449 ( .INP(n2186), .ZN(n2184) );
  INVX0 U2450 ( .INP(n2187), .ZN(n2185) );
  INVX0 U2451 ( .INP(n2190), .ZN(n2188) );
  INVX0 U2452 ( .INP(n2191), .ZN(n2189) );
  INVX0 U2453 ( .INP(n2194), .ZN(n2192) );
  INVX0 U2454 ( .INP(n2195), .ZN(n2193) );
  INVX0 U2455 ( .INP(n2198), .ZN(n2196) );
  INVX0 U2456 ( .INP(n2199), .ZN(n2197) );
  INVX0 U2457 ( .INP(n2202), .ZN(n2200) );
  INVX0 U2458 ( .INP(n2203), .ZN(n2201) );
endmodule


module alu_DW01_add_0 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1, n2;
  wire   [32:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  NAND2X1 U1 ( .IN1(n1), .IN2(n2), .QN(carry[1]) );
  INVX0 U2 ( .INP(A[0]), .ZN(n1) );
  INVX0 U3 ( .INP(B[0]), .ZN(n2) );
  XOR2X1 U4 ( .IN1(n2), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module alu_DW01_add_1 ( A, B, CI, SUM, CO );
  input [32:0] A;
  input [32:0] B;
  output [32:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [32:1] carry;

  FADDX1 U1_31 ( .A(A[31]), .B(B[31]), .CI(carry[31]), .CO(SUM[32]), .S(
        SUM[31]) );
  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  AND2X1 U1 ( .IN1(A[0]), .IN2(B[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[0]), .IN2(B[0]), .Q(SUM[0]) );
endmodule


module alu ( opA, opB, sel, res, z, neg );
  input [31:0] opA;
  input [31:0] opB;
  input [1:0] sel;
  output [31:0] res;
  output z, neg;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N69, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93,
         N94, N95, N96, N97, N98, N99, N100, N101, n10, n11, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n2, n4, n5, n6, n7, n8, n9, n12,
         n13, n24, n25;
  wire   [31:0] res_add;
  wire   [31:0] res_sub;
  assign neg = N101;

  LATCHX1 \res_reg[31]  ( .CLK(n2), .D(N100), .Q(res[31]) );
  LATCHX1 \res_reg[30]  ( .CLK(n2), .D(N99), .Q(res[30]) );
  LATCHX1 \res_reg[29]  ( .CLK(n2), .D(N98), .Q(res[29]) );
  LATCHX1 \res_reg[28]  ( .CLK(n2), .D(N97), .Q(res[28]) );
  LATCHX1 \res_reg[27]  ( .CLK(n2), .D(N96), .Q(res[27]) );
  LATCHX1 \res_reg[26]  ( .CLK(n2), .D(N95), .Q(res[26]) );
  LATCHX1 \res_reg[25]  ( .CLK(n2), .D(N94), .Q(res[25]) );
  LATCHX1 \res_reg[24]  ( .CLK(n2), .D(N93), .Q(res[24]) );
  LATCHX1 \res_reg[23]  ( .CLK(n2), .D(N92), .Q(res[23]) );
  LATCHX1 \res_reg[22]  ( .CLK(n2), .D(N91), .Q(res[22]) );
  LATCHX1 \res_reg[21]  ( .CLK(n2), .D(N90), .Q(res[21]) );
  LATCHX1 \res_reg[20]  ( .CLK(n2), .D(N89), .Q(res[20]) );
  LATCHX1 \res_reg[19]  ( .CLK(n4), .D(N88), .Q(res[19]) );
  LATCHX1 \res_reg[18]  ( .CLK(n4), .D(N87), .Q(res[18]) );
  LATCHX1 \res_reg[17]  ( .CLK(n4), .D(N86), .Q(res[17]) );
  LATCHX1 \res_reg[16]  ( .CLK(n4), .D(N85), .Q(res[16]) );
  LATCHX1 \res_reg[15]  ( .CLK(n4), .D(N84), .Q(res[15]) );
  LATCHX1 \res_reg[14]  ( .CLK(n4), .D(N83), .Q(res[14]) );
  LATCHX1 \res_reg[13]  ( .CLK(n4), .D(N82), .Q(res[13]) );
  LATCHX1 \res_reg[12]  ( .CLK(n4), .D(N81), .Q(res[12]) );
  LATCHX1 \res_reg[11]  ( .CLK(n4), .D(N80), .Q(res[11]) );
  LATCHX1 \res_reg[10]  ( .CLK(n4), .D(N79), .Q(res[10]) );
  LATCHX1 \res_reg[9]  ( .CLK(n4), .D(N78), .Q(res[9]) );
  LATCHX1 \res_reg[8]  ( .CLK(n4), .D(N77), .Q(res[8]) );
  LATCHX1 \res_reg[7]  ( .CLK(n5), .D(N76), .Q(res[7]) );
  LATCHX1 \res_reg[6]  ( .CLK(n5), .D(N75), .Q(res[6]) );
  LATCHX1 \res_reg[5]  ( .CLK(n5), .D(N74), .Q(res[5]) );
  LATCHX1 \res_reg[4]  ( .CLK(n5), .D(N73), .Q(res[4]) );
  LATCHX1 \res_reg[3]  ( .CLK(n5), .D(N72), .Q(res[3]) );
  LATCHX1 \res_reg[2]  ( .CLK(n5), .D(N71), .Q(res[2]) );
  LATCHX1 \res_reg[1]  ( .CLK(n5), .D(N70), .Q(res[1]) );
  LATCHX1 \res_reg[0]  ( .CLK(n5), .D(N69), .Q(res[0]) );
  NAND4X0 U9 ( .IN1(n16), .IN2(n17), .IN3(n18), .IN4(n19), .QN(n15) );
  NOR4X0 U10 ( .IN1(res[23]), .IN2(res[22]), .IN3(res[21]), .IN4(res[20]), 
        .QN(n19) );
  NOR4X0 U11 ( .IN1(res[1]), .IN2(res[19]), .IN3(res[18]), .IN4(res[17]), .QN(
        n18) );
  NOR4X0 U12 ( .IN1(res[16]), .IN2(res[15]), .IN3(res[14]), .IN4(res[13]), 
        .QN(n17) );
  NOR4X0 U13 ( .IN1(res[12]), .IN2(res[11]), .IN3(res[10]), .IN4(res[0]), .QN(
        n16) );
  NAND4X0 U14 ( .IN1(n20), .IN2(n21), .IN3(n22), .IN4(n23), .QN(n14) );
  NOR4X0 U15 ( .IN1(res[9]), .IN2(res[8]), .IN3(res[7]), .IN4(res[6]), .QN(n23) );
  NOR4X0 U16 ( .IN1(res[5]), .IN2(res[4]), .IN3(res[3]), .IN4(res[31]), .QN(
        n22) );
  NOR4X0 U17 ( .IN1(res[30]), .IN2(res[2]), .IN3(res[29]), .IN4(res[28]), .QN(
        n21) );
  NOR4X0 U18 ( .IN1(res[27]), .IN2(res[26]), .IN3(res[25]), .IN4(res[24]), 
        .QN(n20) );
  AO22X1 U19 ( .IN1(n8), .IN2(res_sub[30]), .IN3(res_add[30]), .IN4(n6), .Q(
        N99) );
  AO22X1 U20 ( .IN1(res_sub[29]), .IN2(n8), .IN3(res_add[29]), .IN4(n6), .Q(
        N98) );
  AO22X1 U21 ( .IN1(res_sub[28]), .IN2(n8), .IN3(res_add[28]), .IN4(n6), .Q(
        N97) );
  AO22X1 U22 ( .IN1(res_sub[27]), .IN2(n8), .IN3(res_add[27]), .IN4(n6), .Q(
        N96) );
  AO22X1 U23 ( .IN1(res_sub[26]), .IN2(n9), .IN3(res_add[26]), .IN4(n6), .Q(
        N95) );
  AO22X1 U24 ( .IN1(res_sub[25]), .IN2(n9), .IN3(res_add[25]), .IN4(n6), .Q(
        N94) );
  AO22X1 U25 ( .IN1(res_sub[24]), .IN2(n9), .IN3(res_add[24]), .IN4(n6), .Q(
        N93) );
  AO22X1 U26 ( .IN1(res_sub[23]), .IN2(n9), .IN3(res_add[23]), .IN4(n6), .Q(
        N92) );
  AO22X1 U27 ( .IN1(res_sub[22]), .IN2(n9), .IN3(res_add[22]), .IN4(n6), .Q(
        N91) );
  AO22X1 U28 ( .IN1(res_sub[21]), .IN2(n9), .IN3(res_add[21]), .IN4(n6), .Q(
        N90) );
  AO22X1 U29 ( .IN1(res_sub[20]), .IN2(n9), .IN3(res_add[20]), .IN4(n6), .Q(
        N89) );
  AO22X1 U30 ( .IN1(res_sub[19]), .IN2(n12), .IN3(res_add[19]), .IN4(n6), .Q(
        N88) );
  AO22X1 U31 ( .IN1(res_sub[18]), .IN2(n12), .IN3(res_add[18]), .IN4(n7), .Q(
        N87) );
  AO22X1 U32 ( .IN1(res_sub[17]), .IN2(n12), .IN3(res_add[17]), .IN4(n7), .Q(
        N86) );
  AO22X1 U33 ( .IN1(res_sub[16]), .IN2(n12), .IN3(res_add[16]), .IN4(n7), .Q(
        N85) );
  AO22X1 U34 ( .IN1(res_sub[15]), .IN2(n12), .IN3(res_add[15]), .IN4(n7), .Q(
        N84) );
  AO22X1 U35 ( .IN1(res_sub[14]), .IN2(n12), .IN3(res_add[14]), .IN4(n7), .Q(
        N83) );
  AO22X1 U36 ( .IN1(res_sub[13]), .IN2(n12), .IN3(res_add[13]), .IN4(n7), .Q(
        N82) );
  AO22X1 U37 ( .IN1(res_sub[12]), .IN2(n13), .IN3(res_add[12]), .IN4(n7), .Q(
        N81) );
  AO22X1 U38 ( .IN1(res_sub[11]), .IN2(n13), .IN3(res_add[11]), .IN4(n7), .Q(
        N80) );
  AO22X1 U39 ( .IN1(res_sub[10]), .IN2(n13), .IN3(res_add[10]), .IN4(n7), .Q(
        N79) );
  AO22X1 U40 ( .IN1(res_sub[9]), .IN2(n13), .IN3(res_add[9]), .IN4(n7), .Q(N78) );
  AO22X1 U41 ( .IN1(res_sub[8]), .IN2(n13), .IN3(res_add[8]), .IN4(n7), .Q(N77) );
  AO22X1 U42 ( .IN1(res_sub[7]), .IN2(n13), .IN3(res_add[7]), .IN4(n7), .Q(N76) );
  AO22X1 U43 ( .IN1(res_sub[6]), .IN2(n13), .IN3(res_add[6]), .IN4(n7), .Q(N75) );
  AO22X1 U44 ( .IN1(res_sub[5]), .IN2(n24), .IN3(res_add[5]), .IN4(n6), .Q(N74) );
  AO22X1 U45 ( .IN1(res_sub[4]), .IN2(n24), .IN3(res_add[4]), .IN4(n7), .Q(N73) );
  AO22X1 U46 ( .IN1(res_sub[3]), .IN2(n24), .IN3(res_add[3]), .IN4(n6), .Q(N72) );
  AO22X1 U47 ( .IN1(res_sub[2]), .IN2(n24), .IN3(res_add[2]), .IN4(n7), .Q(N71) );
  AO22X1 U48 ( .IN1(res_sub[1]), .IN2(n24), .IN3(res_add[1]), .IN4(n6), .Q(N70) );
  AO22X1 U49 ( .IN1(res_sub[0]), .IN2(n24), .IN3(res_add[0]), .IN4(n7), .Q(N69) );
  AND3X1 U50 ( .IN1(n11), .IN2(n10), .IN3(res_sub[31]), .Q(N101) );
  AO22X1 U51 ( .IN1(res_sub[31]), .IN2(n24), .IN3(res_add[31]), .IN4(n6), .Q(
        N100) );
  alu_DW01_add_0 add_1_root_add_17_2 ( .A({1'b0, opA}), .B({1'b0, N2, N3, N4, 
        N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, 
        N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33}), 
        .CI(1'b1), .SUM({n10, res_sub}) );
  alu_DW01_add_1 add_16 ( .A({1'b0, opA}), .B({1'b0, opB}), .CI(1'b0), .SUM({
        n11, res_add}) );
  INVX0 U3 ( .INP(opB[9]), .ZN(N24) );
  INVX0 U4 ( .INP(opB[10]), .ZN(N23) );
  INVX0 U6 ( .INP(opB[11]), .ZN(N22) );
  INVX0 U8 ( .INP(opB[15]), .ZN(N18) );
  INVX0 U52 ( .INP(opB[16]), .ZN(N17) );
  INVX0 U53 ( .INP(opB[18]), .ZN(N15) );
  INVX0 U54 ( .INP(opB[19]), .ZN(N14) );
  INVX0 U55 ( .INP(opB[20]), .ZN(N13) );
  INVX0 U56 ( .INP(opB[21]), .ZN(N12) );
  INVX0 U57 ( .INP(opB[26]), .ZN(N7) );
  INVX0 U58 ( .INP(opB[27]), .ZN(N6) );
  INVX0 U59 ( .INP(opB[8]), .ZN(N25) );
  INVX0 U60 ( .INP(opB[12]), .ZN(N21) );
  INVX0 U61 ( .INP(opB[13]), .ZN(N20) );
  INVX0 U62 ( .INP(opB[14]), .ZN(N19) );
  INVX0 U63 ( .INP(opB[17]), .ZN(N16) );
  INVX0 U64 ( .INP(opB[22]), .ZN(N11) );
  INVX0 U65 ( .INP(opB[23]), .ZN(N10) );
  INVX0 U66 ( .INP(opB[24]), .ZN(N9) );
  INVX0 U67 ( .INP(opB[25]), .ZN(N8) );
  INVX0 U68 ( .INP(opB[28]), .ZN(N5) );
  INVX0 U69 ( .INP(opB[29]), .ZN(N4) );
  INVX0 U70 ( .INP(opB[30]), .ZN(N3) );
  INVX0 U71 ( .INP(opB[1]), .ZN(N32) );
  INVX0 U72 ( .INP(opB[2]), .ZN(N31) );
  INVX0 U73 ( .INP(opB[3]), .ZN(N30) );
  INVX0 U74 ( .INP(opB[4]), .ZN(N29) );
  INVX0 U75 ( .INP(opB[5]), .ZN(N28) );
  INVX0 U76 ( .INP(opB[6]), .ZN(N27) );
  INVX0 U77 ( .INP(opB[7]), .ZN(N26) );
  INVX0 U78 ( .INP(opB[31]), .ZN(N2) );
  INVX0 U79 ( .INP(opB[0]), .ZN(N33) );
  NBUFFX2 U80 ( .INP(n25), .Z(n4) );
  NBUFFX2 U81 ( .INP(n25), .Z(n2) );
  NBUFFX2 U82 ( .INP(n25), .Z(n5) );
  NBUFFX2 U83 ( .INP(sel[0]), .Z(n8) );
  NBUFFX2 U84 ( .INP(sel[0]), .Z(n13) );
  NBUFFX2 U85 ( .INP(sel[0]), .Z(n12) );
  NBUFFX2 U86 ( .INP(sel[0]), .Z(n9) );
  NBUFFX2 U87 ( .INP(sel[0]), .Z(n24) );
  INVX0 U88 ( .INP(sel[1]), .ZN(n25) );
  NOR2X0 U89 ( .IN1(n14), .IN2(n15), .QN(z) );
  INVX0 U90 ( .INP(n8), .ZN(n6) );
  INVX0 U91 ( .INP(n8), .ZN(n7) );
endmodule


module single_cycle_mips_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [31:1] carry;

  FADDX1 U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  FADDX1 U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  FADDX1 U1_28 ( .A(A[28]), .B(B[28]), .CI(carry[28]), .CO(carry[29]), .S(
        SUM[28]) );
  FADDX1 U1_27 ( .A(A[27]), .B(B[27]), .CI(carry[27]), .CO(carry[28]), .S(
        SUM[27]) );
  FADDX1 U1_26 ( .A(A[26]), .B(B[26]), .CI(carry[26]), .CO(carry[27]), .S(
        SUM[26]) );
  FADDX1 U1_25 ( .A(A[25]), .B(B[25]), .CI(carry[25]), .CO(carry[26]), .S(
        SUM[25]) );
  FADDX1 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  FADDX1 U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(carry[24]), .S(
        SUM[23]) );
  FADDX1 U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1 U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(n1), .CO(carry[4]), .S(SUM[3]) );
  XOR3X1 U1_31 ( .IN1(A[31]), .IN2(B[31]), .IN3(carry[31]), .Q(SUM[31]) );
  AND2X1 U1 ( .IN1(A[2]), .IN2(B[2]), .Q(n1) );
  XOR2X1 U2 ( .IN1(A[2]), .IN2(B[2]), .Q(SUM[2]) );
endmodule


module single_cycle_mips_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28;

  AND2X1 U1 ( .IN1(A[30]), .IN2(n28), .Q(n1) );
  AND2X1 U2 ( .IN1(A[4]), .IN2(n19), .Q(n2) );
  AND2X1 U3 ( .IN1(A[5]), .IN2(n2), .Q(n3) );
  AND2X1 U4 ( .IN1(A[6]), .IN2(n3), .Q(n4) );
  AND2X1 U5 ( .IN1(A[7]), .IN2(n4), .Q(n5) );
  AND2X1 U6 ( .IN1(A[8]), .IN2(n5), .Q(n6) );
  AND2X1 U7 ( .IN1(A[9]), .IN2(n6), .Q(n7) );
  AND2X1 U8 ( .IN1(A[10]), .IN2(n7), .Q(n8) );
  AND2X1 U9 ( .IN1(A[12]), .IN2(n20), .Q(n9) );
  AND2X1 U10 ( .IN1(A[13]), .IN2(n9), .Q(n10) );
  AND2X1 U11 ( .IN1(A[14]), .IN2(n10), .Q(n11) );
  AND2X1 U12 ( .IN1(A[16]), .IN2(n21), .Q(n12) );
  AND2X1 U13 ( .IN1(A[17]), .IN2(n12), .Q(n13) );
  AND2X1 U14 ( .IN1(A[18]), .IN2(n13), .Q(n14) );
  AND2X1 U15 ( .IN1(A[19]), .IN2(n14), .Q(n15) );
  AND2X1 U16 ( .IN1(A[20]), .IN2(n15), .Q(n16) );
  AND2X1 U17 ( .IN1(A[21]), .IN2(n16), .Q(n17) );
  AND2X1 U18 ( .IN1(A[22]), .IN2(n17), .Q(n18) );
  AND2X1 U19 ( .IN1(A[3]), .IN2(A[2]), .Q(n19) );
  AND2X1 U20 ( .IN1(A[11]), .IN2(n8), .Q(n20) );
  AND2X1 U21 ( .IN1(A[15]), .IN2(n11), .Q(n21) );
  AND2X1 U22 ( .IN1(A[23]), .IN2(n18), .Q(n22) );
  AND2X1 U23 ( .IN1(A[24]), .IN2(n22), .Q(n23) );
  AND2X1 U24 ( .IN1(A[25]), .IN2(n23), .Q(n24) );
  AND2X1 U25 ( .IN1(A[26]), .IN2(n24), .Q(n25) );
  AND2X1 U26 ( .IN1(A[27]), .IN2(n25), .Q(n26) );
  AND2X1 U27 ( .IN1(A[28]), .IN2(n26), .Q(n27) );
  AND2X1 U28 ( .IN1(A[29]), .IN2(n27), .Q(n28) );
  INVX0 U29 ( .INP(A[2]), .ZN(SUM[2]) );
  XOR2X1 U30 ( .IN1(A[31]), .IN2(n1), .Q(SUM[31]) );
  XOR2X1 U31 ( .IN1(A[30]), .IN2(n28), .Q(SUM[30]) );
  XOR2X1 U32 ( .IN1(A[29]), .IN2(n27), .Q(SUM[29]) );
  XOR2X1 U33 ( .IN1(A[28]), .IN2(n26), .Q(SUM[28]) );
  XOR2X1 U34 ( .IN1(A[27]), .IN2(n25), .Q(SUM[27]) );
  XOR2X1 U35 ( .IN1(A[26]), .IN2(n24), .Q(SUM[26]) );
  XOR2X1 U36 ( .IN1(A[25]), .IN2(n23), .Q(SUM[25]) );
  XOR2X1 U37 ( .IN1(A[24]), .IN2(n22), .Q(SUM[24]) );
  XOR2X1 U38 ( .IN1(A[23]), .IN2(n18), .Q(SUM[23]) );
  XOR2X1 U39 ( .IN1(A[22]), .IN2(n17), .Q(SUM[22]) );
  XOR2X1 U40 ( .IN1(A[21]), .IN2(n16), .Q(SUM[21]) );
  XOR2X1 U41 ( .IN1(A[20]), .IN2(n15), .Q(SUM[20]) );
  XOR2X1 U42 ( .IN1(A[19]), .IN2(n14), .Q(SUM[19]) );
  XOR2X1 U43 ( .IN1(A[18]), .IN2(n13), .Q(SUM[18]) );
  XOR2X1 U44 ( .IN1(A[17]), .IN2(n12), .Q(SUM[17]) );
  XOR2X1 U45 ( .IN1(A[16]), .IN2(n21), .Q(SUM[16]) );
  XOR2X1 U46 ( .IN1(A[15]), .IN2(n11), .Q(SUM[15]) );
  XOR2X1 U47 ( .IN1(A[14]), .IN2(n10), .Q(SUM[14]) );
  XOR2X1 U48 ( .IN1(A[13]), .IN2(n9), .Q(SUM[13]) );
  XOR2X1 U49 ( .IN1(A[12]), .IN2(n20), .Q(SUM[12]) );
  XOR2X1 U50 ( .IN1(A[11]), .IN2(n8), .Q(SUM[11]) );
  XOR2X1 U51 ( .IN1(A[10]), .IN2(n7), .Q(SUM[10]) );
  XOR2X1 U52 ( .IN1(A[9]), .IN2(n6), .Q(SUM[9]) );
  XOR2X1 U53 ( .IN1(A[8]), .IN2(n5), .Q(SUM[8]) );
  XOR2X1 U54 ( .IN1(A[7]), .IN2(n4), .Q(SUM[7]) );
  XOR2X1 U55 ( .IN1(A[6]), .IN2(n3), .Q(SUM[6]) );
  XOR2X1 U56 ( .IN1(A[5]), .IN2(n2), .Q(SUM[5]) );
  XOR2X1 U57 ( .IN1(A[4]), .IN2(n19), .Q(SUM[4]) );
  XOR2X1 U58 ( .IN1(A[3]), .IN2(A[2]), .Q(SUM[3]) );
endmodule


module single_cycle_mips ( clk, rst_n, inst_addr, inst, data_addr, data_in, 
        data_out, data_wr );
  output [31:0] inst_addr;
  input [31:0] inst;
  output [31:0] data_addr;
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, rst_n;
  output data_wr;
  wire   aluZ, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66,
         N67, N68, N69, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N460, N461, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88;
  wire   [31:0] rd_dataA;
  wire   [4:0] wr_addr;
  wire   [31:0] wr_data;
  wire   [31:0] aluOpB;
  wire   [1:0] aluSel;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3;
  assign inst_addr[1] = 1'b0;
  assign inst_addr[0] = 1'b0;

  LATCHX1 \aluSel_reg[0]  ( .CLK(N461), .D(N460), .Q(aluSel[0]) );
  LATCHX1 \wr_data_reg[0]  ( .CLK(n55), .D(N522), .Q(wr_data[0]) );
  DFFARX1 \inst_addr_reg[2]  ( .D(N329), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[2]) );
  DFFARX1 \inst_addr_reg[3]  ( .D(N330), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[3]) );
  DFFARX1 \inst_addr_reg[4]  ( .D(N331), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[4]) );
  DFFARX1 \inst_addr_reg[5]  ( .D(N332), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[5]) );
  DFFARX1 \inst_addr_reg[6]  ( .D(N333), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[6]) );
  DFFARX1 \inst_addr_reg[7]  ( .D(N334), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[7]) );
  DFFARX1 \inst_addr_reg[8]  ( .D(N335), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[8]) );
  DFFARX1 \inst_addr_reg[9]  ( .D(N336), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[9]) );
  DFFARX1 \inst_addr_reg[10]  ( .D(N337), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[10]) );
  DFFARX1 \inst_addr_reg[11]  ( .D(N338), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[11]) );
  DFFARX1 \inst_addr_reg[12]  ( .D(N339), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[12]) );
  DFFARX1 \inst_addr_reg[13]  ( .D(N340), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[13]) );
  DFFARX1 \inst_addr_reg[14]  ( .D(N341), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[14]) );
  DFFARX1 \inst_addr_reg[15]  ( .D(N342), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[15]) );
  DFFARX1 \inst_addr_reg[16]  ( .D(N343), .CLK(clk), .RSTB(n74), .Q(
        inst_addr[16]) );
  DFFARX1 \inst_addr_reg[17]  ( .D(N344), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[17]) );
  DFFARX1 \inst_addr_reg[18]  ( .D(N345), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[18]) );
  DFFARX1 \inst_addr_reg[19]  ( .D(N346), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[19]) );
  DFFARX1 \inst_addr_reg[20]  ( .D(N347), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[20]) );
  DFFARX1 \inst_addr_reg[21]  ( .D(N348), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[21]) );
  DFFARX1 \inst_addr_reg[22]  ( .D(N349), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[22]) );
  DFFARX1 \inst_addr_reg[23]  ( .D(N350), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[23]) );
  DFFARX1 \inst_addr_reg[24]  ( .D(N351), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[24]) );
  DFFARX1 \inst_addr_reg[25]  ( .D(N352), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[25]) );
  DFFARX1 \inst_addr_reg[26]  ( .D(N353), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[26]) );
  DFFARX1 \inst_addr_reg[27]  ( .D(N354), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[27]) );
  DFFARX1 \inst_addr_reg[28]  ( .D(N355), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[28]) );
  DFFARX1 \inst_addr_reg[29]  ( .D(N356), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[29]) );
  DFFARX1 \inst_addr_reg[30]  ( .D(N357), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[30]) );
  DFFARX1 \inst_addr_reg[31]  ( .D(N358), .CLK(clk), .RSTB(n56), .Q(
        inst_addr[31]) );
  LATCHX1 \wr_data_reg[1]  ( .CLK(n55), .D(N523), .Q(wr_data[1]) );
  LATCHX1 \wr_data_reg[2]  ( .CLK(n55), .D(N524), .Q(wr_data[2]) );
  LATCHX1 \wr_data_reg[3]  ( .CLK(n55), .D(N525), .Q(wr_data[3]) );
  LATCHX1 \wr_data_reg[4]  ( .CLK(n55), .D(N526), .Q(wr_data[4]) );
  LATCHX1 \wr_data_reg[5]  ( .CLK(n55), .D(N527), .Q(wr_data[5]) );
  LATCHX1 \wr_data_reg[6]  ( .CLK(n55), .D(N528), .Q(wr_data[6]) );
  LATCHX1 \wr_data_reg[7]  ( .CLK(n55), .D(N529), .Q(wr_data[7]) );
  LATCHX1 \wr_data_reg[8]  ( .CLK(n55), .D(N530), .Q(wr_data[8]) );
  LATCHX1 \wr_data_reg[9]  ( .CLK(n55), .D(N531), .Q(wr_data[9]) );
  LATCHX1 \wr_data_reg[10]  ( .CLK(n55), .D(N532), .Q(wr_data[10]) );
  LATCHX1 \wr_data_reg[11]  ( .CLK(n55), .D(N533), .Q(wr_data[11]) );
  LATCHX1 \wr_data_reg[12]  ( .CLK(n55), .D(N534), .Q(wr_data[12]) );
  LATCHX1 \wr_data_reg[13]  ( .CLK(n55), .D(N535), .Q(wr_data[13]) );
  LATCHX1 \wr_data_reg[14]  ( .CLK(n55), .D(N536), .Q(wr_data[14]) );
  LATCHX1 \wr_data_reg[15]  ( .CLK(n55), .D(N537), .Q(wr_data[15]) );
  LATCHX1 \wr_data_reg[16]  ( .CLK(n55), .D(N538), .Q(wr_data[16]) );
  LATCHX1 \wr_data_reg[17]  ( .CLK(n55), .D(N539), .Q(wr_data[17]) );
  LATCHX1 \wr_data_reg[18]  ( .CLK(n55), .D(N540), .Q(wr_data[18]) );
  LATCHX1 \wr_data_reg[19]  ( .CLK(n55), .D(N541), .Q(wr_data[19]) );
  LATCHX1 \wr_data_reg[20]  ( .CLK(n55), .D(N542), .Q(wr_data[20]) );
  LATCHX1 \wr_data_reg[21]  ( .CLK(n55), .D(N543), .Q(wr_data[21]) );
  LATCHX1 \wr_data_reg[22]  ( .CLK(n55), .D(N544), .Q(wr_data[22]) );
  LATCHX1 \wr_data_reg[23]  ( .CLK(n55), .D(N545), .Q(wr_data[23]) );
  LATCHX1 \wr_data_reg[24]  ( .CLK(n55), .D(N546), .Q(wr_data[24]) );
  LATCHX1 \wr_data_reg[25]  ( .CLK(n55), .D(N547), .Q(wr_data[25]) );
  LATCHX1 \wr_data_reg[26]  ( .CLK(n55), .D(N548), .Q(wr_data[26]) );
  LATCHX1 \wr_data_reg[27]  ( .CLK(n55), .D(N549), .Q(wr_data[27]) );
  LATCHX1 \wr_data_reg[28]  ( .CLK(n55), .D(N550), .Q(wr_data[28]) );
  LATCHX1 \wr_data_reg[29]  ( .CLK(n55), .D(N551), .Q(wr_data[29]) );
  LATCHX1 \wr_data_reg[30]  ( .CLK(n55), .D(N552), .Q(wr_data[30]) );
  LATCHX1 \wr_data_reg[31]  ( .CLK(n55), .D(N553), .Q(wr_data[31]) );
  AO22X1 U32 ( .IN1(inst[15]), .IN2(n71), .IN3(inst[20]), .IN4(n25), .Q(
        wr_addr[4]) );
  AO22X1 U33 ( .IN1(inst[14]), .IN2(n72), .IN3(inst[19]), .IN4(n58), .Q(
        wr_addr[3]) );
  AO22X1 U34 ( .IN1(inst[13]), .IN2(n72), .IN3(inst[18]), .IN4(n57), .Q(
        wr_addr[2]) );
  AO22X1 U35 ( .IN1(inst[12]), .IN2(n72), .IN3(inst[17]), .IN4(n25), .Q(
        wr_addr[1]) );
  AO22X1 U36 ( .IN1(inst[11]), .IN2(n72), .IN3(inst[16]), .IN4(n58), .Q(
        wr_addr[0]) );
  AND3X1 U37 ( .IN1(n26), .IN2(inst[29]), .IN3(n83), .Q(data_wr) );
  AO22X1 U38 ( .IN1(data_out[9]), .IN2(n72), .IN3(inst[9]), .IN4(n57), .Q(
        aluOpB[9]) );
  AO22X1 U39 ( .IN1(data_out[8]), .IN2(n72), .IN3(inst[8]), .IN4(n25), .Q(
        aluOpB[8]) );
  AO22X1 U40 ( .IN1(data_out[7]), .IN2(n72), .IN3(inst[7]), .IN4(n58), .Q(
        aluOpB[7]) );
  AO22X1 U41 ( .IN1(data_out[6]), .IN2(n72), .IN3(inst[6]), .IN4(n57), .Q(
        aluOpB[6]) );
  AO22X1 U42 ( .IN1(data_out[5]), .IN2(n72), .IN3(inst[5]), .IN4(n25), .Q(
        aluOpB[5]) );
  AO22X1 U43 ( .IN1(data_out[4]), .IN2(n72), .IN3(inst[4]), .IN4(n58), .Q(
        aluOpB[4]) );
  AO22X1 U44 ( .IN1(data_out[3]), .IN2(n72), .IN3(inst[3]), .IN4(n57), .Q(
        aluOpB[3]) );
  AO21X1 U45 ( .IN1(data_out[31]), .IN2(n70), .IN3(n27), .Q(aluOpB[31]) );
  AO21X1 U46 ( .IN1(data_out[30]), .IN2(n70), .IN3(n27), .Q(aluOpB[30]) );
  AO22X1 U47 ( .IN1(data_out[2]), .IN2(n72), .IN3(inst[2]), .IN4(n25), .Q(
        aluOpB[2]) );
  AO21X1 U48 ( .IN1(data_out[29]), .IN2(n70), .IN3(n27), .Q(aluOpB[29]) );
  AO21X1 U49 ( .IN1(data_out[28]), .IN2(n70), .IN3(n27), .Q(aluOpB[28]) );
  AO21X1 U50 ( .IN1(data_out[27]), .IN2(n71), .IN3(n27), .Q(aluOpB[27]) );
  AO21X1 U51 ( .IN1(data_out[26]), .IN2(n71), .IN3(n27), .Q(aluOpB[26]) );
  AO21X1 U52 ( .IN1(data_out[25]), .IN2(n70), .IN3(n27), .Q(aluOpB[25]) );
  AO21X1 U53 ( .IN1(data_out[24]), .IN2(n71), .IN3(n27), .Q(aluOpB[24]) );
  AO21X1 U54 ( .IN1(data_out[23]), .IN2(n71), .IN3(n27), .Q(aluOpB[23]) );
  AO21X1 U55 ( .IN1(data_out[22]), .IN2(n71), .IN3(n27), .Q(aluOpB[22]) );
  AO21X1 U56 ( .IN1(data_out[21]), .IN2(n70), .IN3(n27), .Q(aluOpB[21]) );
  AO21X1 U57 ( .IN1(data_out[20]), .IN2(n70), .IN3(n27), .Q(aluOpB[20]) );
  AO22X1 U58 ( .IN1(data_out[1]), .IN2(n71), .IN3(inst[1]), .IN4(n58), .Q(
        aluOpB[1]) );
  AO21X1 U59 ( .IN1(data_out[19]), .IN2(n70), .IN3(n27), .Q(aluOpB[19]) );
  AO21X1 U60 ( .IN1(data_out[18]), .IN2(n70), .IN3(n27), .Q(aluOpB[18]) );
  AO21X1 U61 ( .IN1(data_out[17]), .IN2(n70), .IN3(n27), .Q(aluOpB[17]) );
  AO21X1 U62 ( .IN1(data_out[16]), .IN2(n70), .IN3(n27), .Q(aluOpB[16]) );
  AO21X1 U63 ( .IN1(data_out[15]), .IN2(n70), .IN3(n27), .Q(aluOpB[15]) );
  AO22X1 U65 ( .IN1(data_out[14]), .IN2(n71), .IN3(inst[14]), .IN4(n57), .Q(
        aluOpB[14]) );
  AO22X1 U66 ( .IN1(data_out[13]), .IN2(n71), .IN3(inst[13]), .IN4(n25), .Q(
        aluOpB[13]) );
  AO22X1 U67 ( .IN1(data_out[12]), .IN2(n71), .IN3(inst[12]), .IN4(n58), .Q(
        aluOpB[12]) );
  AO22X1 U68 ( .IN1(data_out[11]), .IN2(n71), .IN3(inst[11]), .IN4(n57), .Q(
        aluOpB[11]) );
  AO22X1 U69 ( .IN1(data_out[10]), .IN2(n71), .IN3(inst[10]), .IN4(n25), .Q(
        aluOpB[10]) );
  AO22X1 U70 ( .IN1(data_out[0]), .IN2(n71), .IN3(inst[0]), .IN4(n58), .Q(
        aluOpB[0]) );
  AO221X1 U71 ( .IN1(n29), .IN2(n86), .IN3(inst[26]), .IN4(n30), .IN5(n31), 
        .Q(n24) );
  AO22X1 U73 ( .IN1(data_in[31]), .IN2(n68), .IN3(data_addr[31]), .IN4(n65), 
        .Q(N553) );
  AO22X1 U74 ( .IN1(data_in[30]), .IN2(n69), .IN3(data_addr[30]), .IN4(n65), 
        .Q(N552) );
  AO22X1 U75 ( .IN1(data_in[29]), .IN2(n69), .IN3(data_addr[29]), .IN4(n65), 
        .Q(N551) );
  AO22X1 U76 ( .IN1(data_in[28]), .IN2(n69), .IN3(data_addr[28]), .IN4(n65), 
        .Q(N550) );
  AO22X1 U77 ( .IN1(data_in[27]), .IN2(n69), .IN3(data_addr[27]), .IN4(n65), 
        .Q(N549) );
  AO22X1 U78 ( .IN1(data_in[26]), .IN2(n69), .IN3(data_addr[26]), .IN4(n65), 
        .Q(N548) );
  AO22X1 U79 ( .IN1(data_in[25]), .IN2(n69), .IN3(data_addr[25]), .IN4(n65), 
        .Q(N547) );
  AO22X1 U80 ( .IN1(data_in[24]), .IN2(n69), .IN3(data_addr[24]), .IN4(n65), 
        .Q(N546) );
  AO22X1 U81 ( .IN1(data_in[23]), .IN2(n69), .IN3(data_addr[23]), .IN4(n65), 
        .Q(N545) );
  AO22X1 U82 ( .IN1(data_in[22]), .IN2(n69), .IN3(data_addr[22]), .IN4(n65), 
        .Q(N544) );
  AO22X1 U83 ( .IN1(data_in[21]), .IN2(n69), .IN3(data_addr[21]), .IN4(n65), 
        .Q(N543) );
  AO22X1 U84 ( .IN1(data_in[20]), .IN2(n69), .IN3(data_addr[20]), .IN4(n65), 
        .Q(N542) );
  AO22X1 U85 ( .IN1(data_in[19]), .IN2(n69), .IN3(data_addr[19]), .IN4(n66), 
        .Q(N541) );
  AO22X1 U86 ( .IN1(data_in[18]), .IN2(n68), .IN3(data_addr[18]), .IN4(n66), 
        .Q(N540) );
  AO22X1 U87 ( .IN1(data_in[17]), .IN2(n68), .IN3(data_addr[17]), .IN4(n66), 
        .Q(N539) );
  AO22X1 U88 ( .IN1(data_in[16]), .IN2(n68), .IN3(data_addr[16]), .IN4(n66), 
        .Q(N538) );
  AO22X1 U89 ( .IN1(data_in[15]), .IN2(n68), .IN3(data_addr[15]), .IN4(n66), 
        .Q(N537) );
  AO22X1 U90 ( .IN1(data_in[14]), .IN2(n68), .IN3(data_addr[14]), .IN4(n66), 
        .Q(N536) );
  AO22X1 U91 ( .IN1(data_in[13]), .IN2(n68), .IN3(data_addr[13]), .IN4(n66), 
        .Q(N535) );
  AO22X1 U92 ( .IN1(data_in[12]), .IN2(n68), .IN3(data_addr[12]), .IN4(n66), 
        .Q(N534) );
  AO22X1 U93 ( .IN1(data_in[11]), .IN2(n68), .IN3(data_addr[11]), .IN4(n66), 
        .Q(N533) );
  AO22X1 U94 ( .IN1(data_in[10]), .IN2(n68), .IN3(data_addr[10]), .IN4(n66), 
        .Q(N532) );
  AO22X1 U95 ( .IN1(data_in[9]), .IN2(n68), .IN3(data_addr[9]), .IN4(n66), .Q(
        N531) );
  AO22X1 U96 ( .IN1(data_in[8]), .IN2(n68), .IN3(data_addr[8]), .IN4(n66), .Q(
        N530) );
  AO22X1 U97 ( .IN1(data_in[7]), .IN2(n68), .IN3(data_addr[7]), .IN4(n67), .Q(
        N529) );
  AO22X1 U98 ( .IN1(data_in[6]), .IN2(n68), .IN3(data_addr[6]), .IN4(n67), .Q(
        N528) );
  AO22X1 U99 ( .IN1(data_in[5]), .IN2(n68), .IN3(data_addr[5]), .IN4(n67), .Q(
        N527) );
  AO22X1 U100 ( .IN1(data_in[4]), .IN2(n68), .IN3(data_addr[4]), .IN4(n67), 
        .Q(N526) );
  AO22X1 U101 ( .IN1(data_in[3]), .IN2(n68), .IN3(data_addr[3]), .IN4(n67), 
        .Q(N525) );
  AO22X1 U102 ( .IN1(data_in[2]), .IN2(n68), .IN3(data_addr[2]), .IN4(n67), 
        .Q(N524) );
  AO22X1 U103 ( .IN1(data_in[1]), .IN2(n68), .IN3(data_addr[1]), .IN4(n67), 
        .Q(N523) );
  AO221X1 U104 ( .IN1(data_in[0]), .IN2(n68), .IN3(n87), .IN4(n32), .IN5(n37), 
        .Q(N522) );
  AO21X1 U105 ( .IN1(data_addr[0]), .IN2(n67), .IN3(n33), .Q(n37) );
  AO21X1 U106 ( .IN1(n32), .IN2(n38), .IN3(n34), .Q(n36) );
  NAND4X0 U107 ( .IN1(inst[3]), .IN2(inst[5]), .IN3(inst[1]), .IN4(n39), .QN(
        n38) );
  NOR3X0 U108 ( .IN1(inst[0]), .IN2(inst[4]), .IN3(inst[2]), .QN(n39) );
  AO22X1 U109 ( .IN1(n40), .IN2(n84), .IN3(n83), .IN4(n41), .Q(N461) );
  NAND3X0 U110 ( .IN1(n76), .IN2(n82), .IN3(n42), .QN(n41) );
  NAND4X0 U111 ( .IN1(n43), .IN2(n44), .IN3(inst[5]), .IN4(n45), .QN(n42) );
  NOR4X0 U112 ( .IN1(inst[4]), .IN2(inst[2]), .IN3(inst[26]), .IN4(inst[0]), 
        .QN(n45) );
  AO21X1 U113 ( .IN1(n32), .IN2(inst[1]), .IN3(n40), .Q(N460) );
  AO22X1 U114 ( .IN1(n33), .IN2(n85), .IN3(n47), .IN4(inst[28]), .Q(n40) );
  AND2X1 U115 ( .IN1(inst[27]), .IN2(n46), .Q(n33) );
  AND3X1 U116 ( .IN1(n86), .IN2(n78), .IN3(inst[29]), .Q(n46) );
  AO22X1 U117 ( .IN1(N69), .IN2(n62), .IN3(N101), .IN4(n60), .Q(N358) );
  AO22X1 U118 ( .IN1(N68), .IN2(n62), .IN3(N100), .IN4(n59), .Q(N357) );
  AO22X1 U119 ( .IN1(N67), .IN2(n62), .IN3(N99), .IN4(n60), .Q(N356) );
  AO22X1 U120 ( .IN1(N66), .IN2(n62), .IN3(N98), .IN4(n60), .Q(N355) );
  AO22X1 U121 ( .IN1(N65), .IN2(n62), .IN3(N97), .IN4(n60), .Q(N354) );
  AO22X1 U122 ( .IN1(N64), .IN2(n62), .IN3(N96), .IN4(n60), .Q(N353) );
  AO22X1 U123 ( .IN1(N63), .IN2(n62), .IN3(N95), .IN4(n60), .Q(N352) );
  AO22X1 U124 ( .IN1(N62), .IN2(n62), .IN3(N94), .IN4(n60), .Q(N351) );
  AO22X1 U125 ( .IN1(N61), .IN2(n62), .IN3(N93), .IN4(n60), .Q(N350) );
  AO22X1 U126 ( .IN1(N60), .IN2(n62), .IN3(N92), .IN4(n60), .Q(N349) );
  AO22X1 U127 ( .IN1(N59), .IN2(n62), .IN3(N91), .IN4(n60), .Q(N348) );
  AO22X1 U128 ( .IN1(N58), .IN2(n62), .IN3(N90), .IN4(n60), .Q(N347) );
  AO22X1 U129 ( .IN1(N57), .IN2(n63), .IN3(N89), .IN4(n59), .Q(N346) );
  AO22X1 U130 ( .IN1(N56), .IN2(n63), .IN3(N88), .IN4(n61), .Q(N345) );
  AO22X1 U131 ( .IN1(N55), .IN2(n63), .IN3(N87), .IN4(n59), .Q(N344) );
  AO22X1 U132 ( .IN1(N54), .IN2(n63), .IN3(N86), .IN4(n61), .Q(N343) );
  AO22X1 U133 ( .IN1(N53), .IN2(n63), .IN3(N85), .IN4(n59), .Q(N342) );
  AO22X1 U134 ( .IN1(N52), .IN2(n63), .IN3(N84), .IN4(n61), .Q(N341) );
  AO22X1 U135 ( .IN1(N51), .IN2(n63), .IN3(N83), .IN4(n59), .Q(N340) );
  AO22X1 U136 ( .IN1(N50), .IN2(n63), .IN3(N82), .IN4(n61), .Q(N339) );
  AO22X1 U137 ( .IN1(N49), .IN2(n63), .IN3(N81), .IN4(n59), .Q(N338) );
  AO22X1 U138 ( .IN1(N48), .IN2(n63), .IN3(N80), .IN4(n61), .Q(N337) );
  AO22X1 U139 ( .IN1(N47), .IN2(n63), .IN3(N79), .IN4(n59), .Q(N336) );
  AO22X1 U140 ( .IN1(N46), .IN2(n63), .IN3(N78), .IN4(n61), .Q(N335) );
  AO22X1 U141 ( .IN1(N45), .IN2(n64), .IN3(N77), .IN4(n61), .Q(N334) );
  AO22X1 U142 ( .IN1(N44), .IN2(n64), .IN3(N76), .IN4(n59), .Q(N333) );
  AO22X1 U143 ( .IN1(N43), .IN2(n64), .IN3(N75), .IN4(n61), .Q(N332) );
  AO22X1 U144 ( .IN1(N42), .IN2(n64), .IN3(N74), .IN4(n59), .Q(N331) );
  AO22X1 U145 ( .IN1(N41), .IN2(n64), .IN3(N73), .IN4(n61), .Q(N330) );
  AO22X1 U146 ( .IN1(N40), .IN2(n64), .IN3(N72), .IN4(n59), .Q(N329) );
  AO222X1 U150 ( .IN1(n50), .IN2(n51), .IN3(aluZ), .IN4(n81), .IN5(n79), .IN6(
        n75), .Q(n48) );
  NAND3X0 U151 ( .IN1(n32), .IN2(n84), .IN3(inst[28]), .QN(n51) );
  NOR3X0 U152 ( .IN1(inst[26]), .IN2(inst[29]), .IN3(n80), .QN(n32) );
  NAND4X0 U153 ( .IN1(inst[28]), .IN2(inst[26]), .IN3(n52), .IN4(n43), .QN(n50) );
  rf R1 ( .clk(clk), .rst_n(n73), .rd_addrA(inst[25:21]), .rd_addrB(
        inst[20:16]), .rd_dataA(rd_dataA), .rd_dataB(data_out), .wr_en(n55), 
        .wr_addr(wr_addr), .wr_data(wr_data) );
  alu A1 ( .opA(rd_dataA), .opB(aluOpB), .sel({1'b0, aluSel[0]}), .res(
        data_addr), .z(aluZ) );
  single_cycle_mips_DW01_add_0 r79 ( .A({N69, N68, N67, N66, N65, N64, N63, 
        N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, 
        N48, N47, N46, N45, N44, N43, N42, N41, N40, 1'b0, 1'b0}), .B({
        inst[15], inst[15], inst[15], inst[15], inst[15], inst[15], inst[15], 
        inst[15], inst[15], inst[15], inst[15], inst[15], inst[15], inst[15], 
        inst[15:0], 1'b0, 1'b0}), .CI(1'b0), .SUM({N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, 
        N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1}) );
  single_cycle_mips_DW01_add_1 r78 ( .A({inst_addr[31:2], 1'b0, 1'b0}), .B({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({N69, 
        N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3}) );
  OA21X1 U155 ( .IN1(n28), .IN2(n32), .IN3(n83), .Q(n55) );
  OA21X1 U156 ( .IN1(n28), .IN2(n26), .IN3(n83), .Q(n57) );
  INVX0 U157 ( .INP(n31), .ZN(n83) );
  NBUFFX2 U158 ( .INP(n36), .Z(n65) );
  NBUFFX2 U159 ( .INP(n36), .Z(n66) );
  NBUFFX2 U160 ( .INP(n36), .Z(n67) );
  NBUFFX2 U161 ( .INP(n35), .Z(n68) );
  NBUFFX2 U162 ( .INP(n24), .Z(n71) );
  NBUFFX2 U163 ( .INP(n24), .Z(n72) );
  NAND2X1 U164 ( .IN1(n85), .IN2(n84), .QN(n31) );
  NBUFFX2 U165 ( .INP(n24), .Z(n70) );
  INVX0 U166 ( .INP(n43), .ZN(n80) );
  INVX0 U167 ( .INP(n51), .ZN(n79) );
  INVX0 U168 ( .INP(n50), .ZN(n81) );
  NBUFFX4 U169 ( .INP(n73), .Z(n56) );
  NBUFFX2 U170 ( .INP(n35), .Z(n69) );
  NOR2X0 U171 ( .IN1(n82), .IN2(inst[29]), .QN(n35) );
  INVX0 U172 ( .INP(inst[26]), .ZN(n86) );
  NAND2X0 U173 ( .IN1(inst[31]), .IN2(inst[27]), .QN(n30) );
  AND2X1 U174 ( .IN1(inst[15]), .IN2(n57), .Q(n27) );
  NOR2X0 U175 ( .IN1(n77), .IN2(inst[27]), .QN(n34) );
  INVX0 U176 ( .INP(n46), .ZN(n77) );
  INVX0 U177 ( .INP(inst[31]), .ZN(n78) );
  NAND2X1 U178 ( .IN1(inst[29]), .IN2(n78), .QN(n29) );
  INVX0 U179 ( .INP(inst[30]), .ZN(n84) );
  INVX0 U180 ( .INP(inst[28]), .ZN(n85) );
  NOR2X0 U181 ( .IN1(inst[27]), .IN2(inst[31]), .QN(n43) );
  NOR2X0 U182 ( .IN1(inst[30]), .IN2(inst[29]), .QN(n52) );
  NBUFFX4 U183 ( .INP(rst_n), .Z(n74) );
  NBUFFX2 U184 ( .INP(rst_n), .Z(n73) );
  INVX0 U185 ( .INP(n38), .ZN(n87) );
  NOR2X0 U186 ( .IN1(inst[29]), .IN2(n80), .QN(n47) );
  INVX0 U187 ( .INP(n34), .ZN(n76) );
  NAND2X1 U188 ( .IN1(inst[3]), .IN2(n88), .QN(n44) );
  INVX0 U189 ( .INP(inst[1]), .ZN(n88) );
  INVX0 U192 ( .INP(n26), .ZN(n82) );
  OR3X2 U193 ( .IN1(n33), .IN2(n34), .IN3(n68), .Q(n28) );
  OA21X1 U194 ( .IN1(n28), .IN2(n26), .IN3(n83), .Q(n58) );
  OA21X1 U195 ( .IN1(n28), .IN2(n26), .IN3(n83), .Q(n25) );
  NOR2X0 U196 ( .IN1(n86), .IN2(n30), .QN(n26) );
  AO22X2 U197 ( .IN1(aluZ), .IN2(n79), .IN3(n81), .IN4(n75), .Q(n49) );
  INVX0 U198 ( .INP(aluZ), .ZN(n75) );
  DELLN1X2 U199 ( .INP(n49), .Z(n59) );
  DELLN1X2 U200 ( .INP(n49), .Z(n60) );
  DELLN1X2 U201 ( .INP(n49), .Z(n61) );
  DELLN1X2 U202 ( .INP(n48), .Z(n62) );
  DELLN1X2 U203 ( .INP(n48), .Z(n63) );
  DELLN1X2 U204 ( .INP(n48), .Z(n64) );
endmodule

